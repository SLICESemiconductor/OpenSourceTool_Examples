* NGSPICE file created from sg13g2_IOPadVss_flat.ext - technology: ihp-sg13g2

.subckt sg13g2_IOPadVss_flat vss vdd iovdd iovss
X0 iovss iovdd.t0 dpantenna l=27.78u w=1.26u
X1 iovss iovdd.t0 dpantenna l=27.78u w=1.26u
X2 iovss.t1 iovss dantenna l=27.78u w=1.26u
X3 iovss.t0 iovss dantenna l=27.78u w=1.26u
R0 iovss.n1020 iovss.n1 21.7649
R1 iovss.n1011 iovss.n4 9.0005
R2 iovss.n10 iovss.n4 9.0005
R3 iovss.n1001 iovss.n4 9.0005
R4 iovss.n1009 iovss.n10 9.0005
R5 iovss.n1008 iovss.n10 9.0005
R6 iovss.n1005 iovss.n10 9.0005
R7 iovss.n1003 iovss.n10 9.0005
R8 iovss.n36 iovss.n10 9.0005
R9 iovss.n919 iovss.n10 9.0005
R10 iovss.n921 iovss.n10 9.0005
R11 iovss.n923 iovss.n10 9.0005
R12 iovss.n925 iovss.n10 9.0005
R13 iovss.n927 iovss.n10 9.0005
R14 iovss.n929 iovss.n10 9.0005
R15 iovss.n931 iovss.n10 9.0005
R16 iovss.n933 iovss.n10 9.0005
R17 iovss.n935 iovss.n10 9.0005
R18 iovss.n937 iovss.n10 9.0005
R19 iovss.n939 iovss.n10 9.0005
R20 iovss.n941 iovss.n10 9.0005
R21 iovss.n943 iovss.n10 9.0005
R22 iovss.n945 iovss.n10 9.0005
R23 iovss.n947 iovss.n10 9.0005
R24 iovss.n949 iovss.n10 9.0005
R25 iovss.n951 iovss.n10 9.0005
R26 iovss.n953 iovss.n10 9.0005
R27 iovss.n955 iovss.n10 9.0005
R28 iovss.n957 iovss.n10 9.0005
R29 iovss.n959 iovss.n10 9.0005
R30 iovss.n961 iovss.n10 9.0005
R31 iovss.n963 iovss.n10 9.0005
R32 iovss.n965 iovss.n10 9.0005
R33 iovss.n967 iovss.n10 9.0005
R34 iovss.n969 iovss.n10 9.0005
R35 iovss.n971 iovss.n10 9.0005
R36 iovss.n973 iovss.n10 9.0005
R37 iovss.n975 iovss.n10 9.0005
R38 iovss.n977 iovss.n10 9.0005
R39 iovss.n979 iovss.n10 9.0005
R40 iovss.n981 iovss.n10 9.0005
R41 iovss.n983 iovss.n10 9.0005
R42 iovss.n985 iovss.n10 9.0005
R43 iovss.n987 iovss.n10 9.0005
R44 iovss.n989 iovss.n10 9.0005
R45 iovss.n991 iovss.n10 9.0005
R46 iovss.n993 iovss.n10 9.0005
R47 iovss.n995 iovss.n10 9.0005
R48 iovss.n997 iovss.n10 9.0005
R49 iovss.n1000 iovss.n10 9.0005
R50 iovss.n1001 iovss.n1000 9.0005
R51 iovss.n1001 iovss.n3 9.0005
R52 iovss.n10 iovss.n3 9.0005
R53 iovss.n747 iovss.n394 9.0005
R54 iovss.n742 iovss.n396 9.0005
R55 iovss.n747 iovss.n396 9.0005
R56 iovss.n742 iovss.n393 9.0005
R57 iovss.n747 iovss.n393 9.0005
R58 iovss.n742 iovss.n398 9.0005
R59 iovss.n747 iovss.n398 9.0005
R60 iovss.n742 iovss.n392 9.0005
R61 iovss.n747 iovss.n392 9.0005
R62 iovss.n742 iovss.n400 9.0005
R63 iovss.n747 iovss.n400 9.0005
R64 iovss.n742 iovss.n391 9.0005
R65 iovss.n747 iovss.n391 9.0005
R66 iovss.n742 iovss.n402 9.0005
R67 iovss.n747 iovss.n402 9.0005
R68 iovss.n742 iovss.n390 9.0005
R69 iovss.n747 iovss.n390 9.0005
R70 iovss.n742 iovss.n404 9.0005
R71 iovss.n747 iovss.n404 9.0005
R72 iovss.n742 iovss.n389 9.0005
R73 iovss.n747 iovss.n389 9.0005
R74 iovss.n742 iovss.n406 9.0005
R75 iovss.n747 iovss.n406 9.0005
R76 iovss.n742 iovss.n388 9.0005
R77 iovss.n747 iovss.n388 9.0005
R78 iovss.n742 iovss.n408 9.0005
R79 iovss.n747 iovss.n408 9.0005
R80 iovss.n742 iovss.n387 9.0005
R81 iovss.n747 iovss.n387 9.0005
R82 iovss.n742 iovss.n410 9.0005
R83 iovss.n747 iovss.n410 9.0005
R84 iovss.n742 iovss.n386 9.0005
R85 iovss.n747 iovss.n386 9.0005
R86 iovss.n742 iovss.n412 9.0005
R87 iovss.n747 iovss.n412 9.0005
R88 iovss.n742 iovss.n385 9.0005
R89 iovss.n747 iovss.n385 9.0005
R90 iovss.n742 iovss.n414 9.0005
R91 iovss.n747 iovss.n414 9.0005
R92 iovss.n742 iovss.n384 9.0005
R93 iovss.n747 iovss.n384 9.0005
R94 iovss.n742 iovss.n416 9.0005
R95 iovss.n747 iovss.n416 9.0005
R96 iovss.n742 iovss.n383 9.0005
R97 iovss.n747 iovss.n383 9.0005
R98 iovss.n742 iovss.n418 9.0005
R99 iovss.n747 iovss.n418 9.0005
R100 iovss.n742 iovss.n382 9.0005
R101 iovss.n747 iovss.n382 9.0005
R102 iovss.n742 iovss.n420 9.0005
R103 iovss.n747 iovss.n420 9.0005
R104 iovss.n742 iovss.n381 9.0005
R105 iovss.n747 iovss.n381 9.0005
R106 iovss.n742 iovss.n422 9.0005
R107 iovss.n747 iovss.n422 9.0005
R108 iovss.n742 iovss.n380 9.0005
R109 iovss.n747 iovss.n380 9.0005
R110 iovss.n742 iovss.n424 9.0005
R111 iovss.n747 iovss.n424 9.0005
R112 iovss.n742 iovss.n379 9.0005
R113 iovss.n747 iovss.n379 9.0005
R114 iovss.n742 iovss.n426 9.0005
R115 iovss.n747 iovss.n426 9.0005
R116 iovss.n742 iovss.n378 9.0005
R117 iovss.n747 iovss.n378 9.0005
R118 iovss.n742 iovss.n428 9.0005
R119 iovss.n747 iovss.n428 9.0005
R120 iovss.n742 iovss.n377 9.0005
R121 iovss.n747 iovss.n377 9.0005
R122 iovss.n742 iovss.n430 9.0005
R123 iovss.n747 iovss.n430 9.0005
R124 iovss.n742 iovss.n376 9.0005
R125 iovss.n747 iovss.n376 9.0005
R126 iovss.n742 iovss.n432 9.0005
R127 iovss.n747 iovss.n432 9.0005
R128 iovss.n742 iovss.n375 9.0005
R129 iovss.n747 iovss.n375 9.0005
R130 iovss.n742 iovss.n434 9.0005
R131 iovss.n747 iovss.n434 9.0005
R132 iovss.n742 iovss.n374 9.0005
R133 iovss.n747 iovss.n374 9.0005
R134 iovss.n742 iovss.n436 9.0005
R135 iovss.n747 iovss.n436 9.0005
R136 iovss.n742 iovss.n373 9.0005
R137 iovss.n747 iovss.n373 9.0005
R138 iovss.n742 iovss.n438 9.0005
R139 iovss.n747 iovss.n438 9.0005
R140 iovss.n742 iovss.n372 9.0005
R141 iovss.n747 iovss.n372 9.0005
R142 iovss.n742 iovss.n440 9.0005
R143 iovss.n747 iovss.n440 9.0005
R144 iovss.n742 iovss.n371 9.0005
R145 iovss.n747 iovss.n371 9.0005
R146 iovss.n742 iovss.n441 9.0005
R147 iovss.n747 iovss.n441 9.0005
R148 iovss.n747 iovss.n746 9.0005
R149 iovss.n746 iovss.n745 9.0005
R150 iovss.n746 iovss.n445 9.0005
R151 iovss.n1018 iovss.n3 9.0005
R152 iovss.n1016 iovss.n3 9.0005
R153 iovss.n5 iovss.n3 9.0005
R154 iovss.n745 iovss.n744 9.0005
R155 iovss.n744 iovss.n445 9.0005
R156 iovss.n1018 iovss.n1017 9.0005
R157 iovss.n1017 iovss.n5 9.0005
R158 iovss.n1017 iovss.n1016 9.0005
R159 iovss.n778 iovss.n777 9.0005
R160 iovss.n777 iovss.n774 9.0005
R161 iovss.n778 iovss.n135 9.0005
R162 iovss.n779 iovss.n160 9.0005
R163 iovss.n781 iovss.n160 9.0005
R164 iovss.n783 iovss.n160 9.0005
R165 iovss.n785 iovss.n160 9.0005
R166 iovss.n787 iovss.n160 9.0005
R167 iovss.n789 iovss.n160 9.0005
R168 iovss.n791 iovss.n160 9.0005
R169 iovss.n793 iovss.n160 9.0005
R170 iovss.n795 iovss.n160 9.0005
R171 iovss.n797 iovss.n160 9.0005
R172 iovss.n799 iovss.n160 9.0005
R173 iovss.n801 iovss.n160 9.0005
R174 iovss.n803 iovss.n160 9.0005
R175 iovss.n805 iovss.n160 9.0005
R176 iovss.n807 iovss.n160 9.0005
R177 iovss.n809 iovss.n160 9.0005
R178 iovss.n811 iovss.n160 9.0005
R179 iovss.n813 iovss.n160 9.0005
R180 iovss.n815 iovss.n160 9.0005
R181 iovss.n817 iovss.n160 9.0005
R182 iovss.n819 iovss.n160 9.0005
R183 iovss.n821 iovss.n160 9.0005
R184 iovss.n823 iovss.n160 9.0005
R185 iovss.n825 iovss.n160 9.0005
R186 iovss.n827 iovss.n160 9.0005
R187 iovss.n829 iovss.n160 9.0005
R188 iovss.n831 iovss.n160 9.0005
R189 iovss.n833 iovss.n160 9.0005
R190 iovss.n835 iovss.n160 9.0005
R191 iovss.n837 iovss.n160 9.0005
R192 iovss.n839 iovss.n160 9.0005
R193 iovss.n841 iovss.n160 9.0005
R194 iovss.n843 iovss.n160 9.0005
R195 iovss.n845 iovss.n160 9.0005
R196 iovss.n847 iovss.n160 9.0005
R197 iovss.n849 iovss.n160 9.0005
R198 iovss.n851 iovss.n160 9.0005
R199 iovss.n853 iovss.n160 9.0005
R200 iovss.n855 iovss.n160 9.0005
R201 iovss.n857 iovss.n160 9.0005
R202 iovss.n859 iovss.n160 9.0005
R203 iovss.n861 iovss.n160 9.0005
R204 iovss.n863 iovss.n160 9.0005
R205 iovss.n865 iovss.n160 9.0005
R206 iovss.n867 iovss.n160 9.0005
R207 iovss.n870 iovss.n160 9.0005
R208 iovss.n771 iovss.n160 9.0005
R209 iovss.n872 iovss.n133 9.0005
R210 iovss.n160 iovss.n133 9.0005
R211 iovss.n886 iovss.n135 9.0005
R212 iovss.n160 iovss.n135 9.0005
R213 iovss.n777 iovss.n160 9.0005
R214 iovss.n774 iovss.n135 9.0005
R215 iovss.n899 iovss.n898 9.0005
R216 iovss.n902 iovss.n103 9.0005
R217 iovss.n902 iovss.n106 9.0005
R218 iovss.n902 iovss.n102 9.0005
R219 iovss.n902 iovss.n108 9.0005
R220 iovss.n902 iovss.n101 9.0005
R221 iovss.n902 iovss.n110 9.0005
R222 iovss.n902 iovss.n100 9.0005
R223 iovss.n902 iovss.n901 9.0005
R224 iovss.n902 iovss.n99 9.0005
R225 iovss.n903 iovss.n96 9.0005
R226 iovss.n903 iovss.n902 9.0005
R227 iovss.n700 iovss.n699 9.0005
R228 iovss.n692 iovss.n460 9.0005
R229 iovss.n699 iovss.n460 9.0005
R230 iovss.n692 iovss.n457 9.0005
R231 iovss.n699 iovss.n457 9.0005
R232 iovss.n692 iovss.n463 9.0005
R233 iovss.n699 iovss.n463 9.0005
R234 iovss.n699 iovss.n456 9.0005
R235 iovss.n692 iovss.n455 9.0005
R236 iovss.n699 iovss.n455 9.0005
R237 iovss.n692 iovss.n467 9.0005
R238 iovss.n699 iovss.n467 9.0005
R239 iovss.n692 iovss.n454 9.0005
R240 iovss.n699 iovss.n454 9.0005
R241 iovss.n699 iovss.n698 9.0005
R242 iovss.n699 iovss.n453 9.0005
R243 iovss.n692 iovss.n95 9.0005
R244 iovss.n699 iovss.n95 9.0005
R245 iovss.n907 iovss.n65 9.0005
R246 iovss.n907 iovss.n906 9.0005
R247 iovss.n906 iovss.n74 9.0005
R248 iovss.n906 iovss.n71 9.0005
R249 iovss.n906 iovss.n77 9.0005
R250 iovss.n906 iovss.n70 9.0005
R251 iovss.n906 iovss.n80 9.0005
R252 iovss.n906 iovss.n69 9.0005
R253 iovss.n906 iovss.n90 9.0005
R254 iovss.n906 iovss.n68 9.0005
R255 iovss.n906 iovss.n93 9.0005
R256 iovss.n906 iovss.n67 9.0005
R257 iovss.n905 iovss.n65 9.0005
R258 iovss.n906 iovss.n905 9.0005
R259 iovss.n1013 iovss.n1012 4.50058
R260 iovss.n1017 iovss.n6 4.50058
R261 iovss.n744 iovss.n370 4.50058
R262 iovss.n746 iovss.n737 4.50058
R263 iovss.n777 iovss.n134 4.50058
R264 iovss.n895 iovss.n117 4.50058
R265 iovss.n700 iovss.n450 4.50058
R266 iovss.n690 iovss.n464 4.50058
R267 iovss.n443 iovss.n442 4.4951
R268 iovss.n1001 iovss.n9 4.49246
R269 iovss.n1011 iovss.n1010 4.49246
R270 iovss.n1001 iovss.n34 4.49246
R271 iovss.n1011 iovss.n33 4.49246
R272 iovss.n1002 iovss.n1001 4.49246
R273 iovss.n1011 iovss.n32 4.49246
R274 iovss.n1001 iovss.n56 4.49246
R275 iovss.n1011 iovss.n31 4.49246
R276 iovss.n1001 iovss.n55 4.49246
R277 iovss.n1011 iovss.n30 4.49246
R278 iovss.n1001 iovss.n54 4.49246
R279 iovss.n1011 iovss.n29 4.49246
R280 iovss.n1001 iovss.n53 4.49246
R281 iovss.n1011 iovss.n28 4.49246
R282 iovss.n1001 iovss.n52 4.49246
R283 iovss.n1011 iovss.n27 4.49246
R284 iovss.n1001 iovss.n51 4.49246
R285 iovss.n1011 iovss.n26 4.49246
R286 iovss.n1001 iovss.n50 4.49246
R287 iovss.n1011 iovss.n25 4.49246
R288 iovss.n1001 iovss.n49 4.49246
R289 iovss.n1011 iovss.n24 4.49246
R290 iovss.n1001 iovss.n48 4.49246
R291 iovss.n1011 iovss.n23 4.49246
R292 iovss.n1001 iovss.n47 4.49246
R293 iovss.n1011 iovss.n22 4.49246
R294 iovss.n1001 iovss.n46 4.49246
R295 iovss.n1011 iovss.n21 4.49246
R296 iovss.n1001 iovss.n45 4.49246
R297 iovss.n1011 iovss.n20 4.49246
R298 iovss.n1001 iovss.n44 4.49246
R299 iovss.n1011 iovss.n19 4.49246
R300 iovss.n1001 iovss.n43 4.49246
R301 iovss.n1011 iovss.n18 4.49246
R302 iovss.n1001 iovss.n42 4.49246
R303 iovss.n1011 iovss.n17 4.49246
R304 iovss.n1001 iovss.n41 4.49246
R305 iovss.n1011 iovss.n16 4.49246
R306 iovss.n1001 iovss.n40 4.49246
R307 iovss.n1011 iovss.n15 4.49246
R308 iovss.n1001 iovss.n39 4.49246
R309 iovss.n1011 iovss.n14 4.49246
R310 iovss.n1001 iovss.n38 4.49246
R311 iovss.n1011 iovss.n13 4.49246
R312 iovss.n1001 iovss.n37 4.49246
R313 iovss.n1011 iovss.n12 4.49246
R314 iovss.n1011 iovss.n7 4.49246
R315 iovss.n743 iovss.n742 4.49246
R316 iovss.n736 iovss.n735 4.49246
R317 iovss.n736 iovss.n734 4.49246
R318 iovss.n736 iovss.n733 4.49246
R319 iovss.n736 iovss.n732 4.49246
R320 iovss.n736 iovss.n731 4.49246
R321 iovss.n736 iovss.n730 4.49246
R322 iovss.n736 iovss.n729 4.49246
R323 iovss.n736 iovss.n728 4.49246
R324 iovss.n736 iovss.n727 4.49246
R325 iovss.n736 iovss.n726 4.49246
R326 iovss.n736 iovss.n725 4.49246
R327 iovss.n736 iovss.n724 4.49246
R328 iovss.n736 iovss.n723 4.49246
R329 iovss.n736 iovss.n722 4.49246
R330 iovss.n736 iovss.n721 4.49246
R331 iovss.n736 iovss.n720 4.49246
R332 iovss.n736 iovss.n719 4.49246
R333 iovss.n736 iovss.n718 4.49246
R334 iovss.n736 iovss.n717 4.49246
R335 iovss.n736 iovss.n716 4.49246
R336 iovss.n736 iovss.n715 4.49246
R337 iovss.n736 iovss.n714 4.49246
R338 iovss.n736 iovss.n713 4.49246
R339 iovss.n736 iovss.n712 4.49246
R340 iovss.n776 iovss.n775 4.49246
R341 iovss.n872 iovss.n748 4.49246
R342 iovss.n886 iovss.n159 4.49246
R343 iovss.n872 iovss.n749 4.49246
R344 iovss.n886 iovss.n158 4.49246
R345 iovss.n872 iovss.n750 4.49246
R346 iovss.n886 iovss.n157 4.49246
R347 iovss.n872 iovss.n751 4.49246
R348 iovss.n886 iovss.n156 4.49246
R349 iovss.n872 iovss.n752 4.49246
R350 iovss.n886 iovss.n155 4.49246
R351 iovss.n872 iovss.n753 4.49246
R352 iovss.n886 iovss.n154 4.49246
R353 iovss.n872 iovss.n754 4.49246
R354 iovss.n886 iovss.n153 4.49246
R355 iovss.n872 iovss.n755 4.49246
R356 iovss.n886 iovss.n152 4.49246
R357 iovss.n872 iovss.n756 4.49246
R358 iovss.n886 iovss.n151 4.49246
R359 iovss.n872 iovss.n757 4.49246
R360 iovss.n886 iovss.n150 4.49246
R361 iovss.n872 iovss.n758 4.49246
R362 iovss.n886 iovss.n149 4.49246
R363 iovss.n872 iovss.n759 4.49246
R364 iovss.n886 iovss.n148 4.49246
R365 iovss.n872 iovss.n760 4.49246
R366 iovss.n886 iovss.n147 4.49246
R367 iovss.n872 iovss.n761 4.49246
R368 iovss.n886 iovss.n146 4.49246
R369 iovss.n872 iovss.n762 4.49246
R370 iovss.n886 iovss.n145 4.49246
R371 iovss.n872 iovss.n763 4.49246
R372 iovss.n886 iovss.n144 4.49246
R373 iovss.n872 iovss.n764 4.49246
R374 iovss.n886 iovss.n143 4.49246
R375 iovss.n872 iovss.n765 4.49246
R376 iovss.n886 iovss.n142 4.49246
R377 iovss.n872 iovss.n766 4.49246
R378 iovss.n886 iovss.n141 4.49246
R379 iovss.n872 iovss.n767 4.49246
R380 iovss.n886 iovss.n140 4.49246
R381 iovss.n872 iovss.n768 4.49246
R382 iovss.n886 iovss.n139 4.49246
R383 iovss.n872 iovss.n769 4.49246
R384 iovss.n886 iovss.n138 4.49246
R385 iovss.n872 iovss.n770 4.49246
R386 iovss.n886 iovss.n137 4.49246
R387 iovss.n872 iovss.n871 4.49246
R388 iovss.n886 iovss.n136 4.49246
R389 iovss.n902 iovss.n104 4.49246
R390 iovss.n118 iovss.n96 4.49246
R391 iovss.n899 iovss.n116 4.49246
R392 iovss.n105 iovss.n96 4.49246
R393 iovss.n899 iovss.n115 4.49246
R394 iovss.n107 iovss.n96 4.49246
R395 iovss.n899 iovss.n114 4.49246
R396 iovss.n109 iovss.n96 4.49246
R397 iovss.n900 iovss.n899 4.49246
R398 iovss.n111 iovss.n96 4.49246
R399 iovss.n899 iovss.n97 4.49246
R400 iovss.n459 iovss.n448 4.49246
R401 iovss.n461 iovss.n448 4.49246
R402 iovss.n692 iovss.n691 4.49246
R403 iovss.n466 iovss.n448 4.49246
R404 iovss.n694 iovss.n448 4.49246
R405 iovss.n693 iovss.n692 4.49246
R406 iovss.n451 iovss.n448 4.49246
R407 iovss.n66 iovss.n64 4.49246
R408 iovss.n73 iovss.n65 4.49246
R409 iovss.n76 iovss.n66 4.49246
R410 iovss.n75 iovss.n65 4.49246
R411 iovss.n79 iovss.n66 4.49246
R412 iovss.n78 iovss.n65 4.49246
R413 iovss.n82 iovss.n66 4.49246
R414 iovss.n81 iovss.n65 4.49246
R415 iovss.n92 iovss.n66 4.49246
R416 iovss.n91 iovss.n65 4.49246
R417 iovss.n94 iovss.n66 4.49246
R418 iovss.n0 iovss.t1 3.07412
R419 iovss.n738 iovss.t0 3.07412
R420 iovss.n456 iovss.n1 3.0079
R421 iovss.n698 iovss.n697 3.00565
R422 iovss.n444 iovss.n394 3.00498
R423 iovss.n914 iovss.n58 3.0005
R424 iovss.n916 iovss.n915 3.0005
R425 iovss.n913 iovss.n60 3.0005
R426 iovss.n912 iovss.n911 3.0005
R427 iovss.n62 iovss.n61 3.0005
R428 iovss.n1015 iovss.n4 3.0005
R429 iovss.n695 iovss.n93 3.0005
R430 iovss.n83 iovss.n68 3.0005
R431 iovss.n90 iovss.n89 3.0005
R432 iovss.n88 iovss.n69 3.0005
R433 iovss.n87 iovss.n80 3.0005
R434 iovss.n86 iovss.n70 3.0005
R435 iovss.n85 iovss.n77 3.0005
R436 iovss.n84 iovss.n71 3.0005
R437 iovss.n74 iovss.n63 3.0005
R438 iovss.n908 iovss.n907 3.0005
R439 iovss.n909 iovss.n62 3.0005
R440 iovss.n911 iovss.n910 3.0005
R441 iovss.n60 iovss.n59 3.0005
R442 iovss.n917 iovss.n916 3.0005
R443 iovss.n918 iovss.n58 3.0005
R444 iovss.n1000 iovss.n999 3.0005
R445 iovss.n998 iovss.n997 3.0005
R446 iovss.n996 iovss.n995 3.0005
R447 iovss.n994 iovss.n993 3.0005
R448 iovss.n992 iovss.n991 3.0005
R449 iovss.n990 iovss.n989 3.0005
R450 iovss.n988 iovss.n987 3.0005
R451 iovss.n986 iovss.n985 3.0005
R452 iovss.n984 iovss.n983 3.0005
R453 iovss.n982 iovss.n981 3.0005
R454 iovss.n980 iovss.n979 3.0005
R455 iovss.n978 iovss.n977 3.0005
R456 iovss.n976 iovss.n975 3.0005
R457 iovss.n974 iovss.n973 3.0005
R458 iovss.n972 iovss.n971 3.0005
R459 iovss.n970 iovss.n969 3.0005
R460 iovss.n968 iovss.n967 3.0005
R461 iovss.n966 iovss.n965 3.0005
R462 iovss.n964 iovss.n963 3.0005
R463 iovss.n962 iovss.n961 3.0005
R464 iovss.n960 iovss.n959 3.0005
R465 iovss.n958 iovss.n957 3.0005
R466 iovss.n956 iovss.n955 3.0005
R467 iovss.n954 iovss.n953 3.0005
R468 iovss.n952 iovss.n951 3.0005
R469 iovss.n950 iovss.n949 3.0005
R470 iovss.n948 iovss.n947 3.0005
R471 iovss.n946 iovss.n945 3.0005
R472 iovss.n944 iovss.n943 3.0005
R473 iovss.n942 iovss.n941 3.0005
R474 iovss.n940 iovss.n939 3.0005
R475 iovss.n938 iovss.n937 3.0005
R476 iovss.n936 iovss.n935 3.0005
R477 iovss.n934 iovss.n933 3.0005
R478 iovss.n932 iovss.n931 3.0005
R479 iovss.n930 iovss.n929 3.0005
R480 iovss.n928 iovss.n927 3.0005
R481 iovss.n926 iovss.n925 3.0005
R482 iovss.n924 iovss.n923 3.0005
R483 iovss.n922 iovss.n921 3.0005
R484 iovss.n920 iovss.n919 3.0005
R485 iovss.n36 iovss.n35 3.0005
R486 iovss.n1004 iovss.n1003 3.0005
R487 iovss.n1006 iovss.n1005 3.0005
R488 iovss.n1008 iovss.n1007 3.0005
R489 iovss.n1009 iovss.n8 3.0005
R490 iovss.n1014 iovss.n1013 3.0005
R491 iovss.n905 iovss.n904 3.0005
R492 iovss.n452 iovss.n67 3.0005
R493 iovss.n904 iovss.n95 3.0005
R494 iovss.n453 iovss.n452 3.0005
R495 iovss.n711 iovss.n710 3.0005
R496 iovss.n708 iovss.n446 3.0005
R497 iovss.n706 iovss.n705 3.0005
R498 iovss.n704 iovss.n447 3.0005
R499 iovss.n703 iovss.n702 3.0005
R500 iovss.n780 iovss.n779 3.0005
R501 iovss.n121 iovss.n101 3.0005
R502 iovss.n122 iovss.n108 3.0005
R503 iovss.n123 iovss.n102 3.0005
R504 iovss.n124 iovss.n106 3.0005
R505 iovss.n125 iovss.n103 3.0005
R506 iovss.n898 iovss.n897 3.0005
R507 iovss.n896 iovss.n895 3.0005
R508 iovss.n894 iovss.n126 3.0005
R509 iovss.n129 iovss.n127 3.0005
R510 iovss.n890 iovss.n130 3.0005
R511 iovss.n889 iovss.n131 3.0005
R512 iovss.n888 iovss.n132 3.0005
R513 iovss.n772 iovss.n133 3.0005
R514 iovss.n773 iovss.n771 3.0005
R515 iovss.n870 iovss.n869 3.0005
R516 iovss.n868 iovss.n867 3.0005
R517 iovss.n866 iovss.n865 3.0005
R518 iovss.n864 iovss.n863 3.0005
R519 iovss.n862 iovss.n861 3.0005
R520 iovss.n860 iovss.n859 3.0005
R521 iovss.n858 iovss.n857 3.0005
R522 iovss.n856 iovss.n855 3.0005
R523 iovss.n854 iovss.n853 3.0005
R524 iovss.n852 iovss.n851 3.0005
R525 iovss.n850 iovss.n849 3.0005
R526 iovss.n848 iovss.n847 3.0005
R527 iovss.n846 iovss.n845 3.0005
R528 iovss.n844 iovss.n843 3.0005
R529 iovss.n842 iovss.n841 3.0005
R530 iovss.n840 iovss.n839 3.0005
R531 iovss.n838 iovss.n837 3.0005
R532 iovss.n836 iovss.n835 3.0005
R533 iovss.n834 iovss.n833 3.0005
R534 iovss.n832 iovss.n831 3.0005
R535 iovss.n830 iovss.n829 3.0005
R536 iovss.n828 iovss.n827 3.0005
R537 iovss.n826 iovss.n825 3.0005
R538 iovss.n824 iovss.n823 3.0005
R539 iovss.n822 iovss.n821 3.0005
R540 iovss.n820 iovss.n819 3.0005
R541 iovss.n818 iovss.n817 3.0005
R542 iovss.n816 iovss.n815 3.0005
R543 iovss.n814 iovss.n813 3.0005
R544 iovss.n812 iovss.n811 3.0005
R545 iovss.n810 iovss.n809 3.0005
R546 iovss.n808 iovss.n807 3.0005
R547 iovss.n806 iovss.n805 3.0005
R548 iovss.n804 iovss.n803 3.0005
R549 iovss.n802 iovss.n801 3.0005
R550 iovss.n800 iovss.n799 3.0005
R551 iovss.n798 iovss.n797 3.0005
R552 iovss.n796 iovss.n795 3.0005
R553 iovss.n794 iovss.n793 3.0005
R554 iovss.n792 iovss.n791 3.0005
R555 iovss.n790 iovss.n789 3.0005
R556 iovss.n788 iovss.n787 3.0005
R557 iovss.n786 iovss.n785 3.0005
R558 iovss.n784 iovss.n783 3.0005
R559 iovss.n782 iovss.n781 3.0005
R560 iovss.n901 iovss.n112 3.0005
R561 iovss.n904 iovss.n903 3.0005
R562 iovss.n452 iovss.n99 3.0005
R563 iovss.n119 iovss.n100 3.0005
R564 iovss.n120 iovss.n110 3.0005
R565 iovss.n888 iovss.n887 3.0005
R566 iovss.n889 iovss.n128 3.0005
R567 iovss.n891 iovss.n890 3.0005
R568 iovss.n892 iovss.n127 3.0005
R569 iovss.n894 iovss.n893 3.0005
R570 iovss.n437 iovss.n1 1.49548
R571 iovss.n403 iovss.n1 1.49548
R572 iovss.n421 iovss.n1 1.49545
R573 iovss.n419 iovss.n1 1.4954
R574 iovss.n439 iovss.n1 1.49532
R575 iovss.n405 iovss.n1 1.49532
R576 iovss.n435 iovss.n1 1.49522
R577 iovss.n401 iovss.n1 1.49522
R578 iovss.n423 iovss.n1 1.49509
R579 iovss.n465 iovss.n1 1.49504
R580 iovss.n429 iovss.n1 1.49504
R581 iovss.n395 iovss.n1 1.49504
R582 iovss.n701 iovss.n1 1.49502
R583 iovss.n411 iovss.n1 1.49502
R584 iovss.n413 iovss.n1 1.49496
R585 iovss.n449 iovss.n1 1.49496
R586 iovss.n417 iovss.n1 1.49494
R587 iovss.n427 iovss.n1 1.49489
R588 iovss.n431 iovss.n1 1.49478
R589 iovss.n397 iovss.n1 1.49478
R590 iovss.n689 iovss.n1 1.49478
R591 iovss.n709 iovss.n1 1.49476
R592 iovss.n407 iovss.n1 1.49476
R593 iovss.n707 iovss.n1 1.49466
R594 iovss.n409 iovss.n1 1.49466
R595 iovss.n433 iovss.n1 1.49455
R596 iovss.n399 iovss.n1 1.49455
R597 iovss.n415 iovss.n1 1.4945
R598 iovss.n462 iovss.n1 1.4945
R599 iovss.n425 iovss.n1 1.49432
R600 iovss.n242 iovss.n239 0.826084
R601 iovss.n546 iovss.n545 0.826084
R602 iovss.n884 iovss.n883 0.822133
R603 iovss.n679 iovss.n678 0.822133
R604 iovss.n241 iovss.n240 0.818682
R605 iovss.n248 iovss.n247 0.818682
R606 iovss.n238 iovss.n236 0.818682
R607 iovss.n253 iovss.n252 0.818682
R608 iovss.n232 iovss.n231 0.818682
R609 iovss.n263 iovss.n262 0.818682
R610 iovss.n229 iovss.n227 0.818682
R611 iovss.n268 iovss.n267 0.818682
R612 iovss.n223 iovss.n222 0.818682
R613 iovss.n278 iovss.n277 0.818682
R614 iovss.n220 iovss.n218 0.818682
R615 iovss.n283 iovss.n282 0.818682
R616 iovss.n214 iovss.n213 0.818682
R617 iovss.n293 iovss.n292 0.818682
R618 iovss.n211 iovss.n209 0.818682
R619 iovss.n298 iovss.n297 0.818682
R620 iovss.n205 iovss.n204 0.818682
R621 iovss.n308 iovss.n307 0.818682
R622 iovss.n202 iovss.n200 0.818682
R623 iovss.n313 iovss.n312 0.818682
R624 iovss.n196 iovss.n195 0.818682
R625 iovss.n323 iovss.n322 0.818682
R626 iovss.n193 iovss.n191 0.818682
R627 iovss.n328 iovss.n327 0.818682
R628 iovss.n187 iovss.n186 0.818682
R629 iovss.n338 iovss.n337 0.818682
R630 iovss.n184 iovss.n182 0.818682
R631 iovss.n343 iovss.n342 0.818682
R632 iovss.n178 iovss.n177 0.818682
R633 iovss.n353 iovss.n352 0.818682
R634 iovss.n175 iovss.n173 0.818682
R635 iovss.n358 iovss.n357 0.818682
R636 iovss.n169 iovss.n168 0.818682
R637 iovss.n368 iovss.n367 0.818682
R638 iovss.n369 iovss.n166 0.818682
R639 iovss.n876 iovss.n875 0.818682
R640 iovss.n162 iovss.n161 0.818682
R641 iovss.n885 iovss.n884 0.818682
R642 iovss.n873 iovss.n161 0.818682
R643 iovss.n875 iovss.n874 0.818682
R644 iovss.n741 iovss.n369 0.818682
R645 iovss.n368 iovss.n57 0.818682
R646 iovss.n168 iovss.n11 0.818682
R647 iovss.n357 iovss.n356 0.818682
R648 iovss.n355 iovss.n175 0.818682
R649 iovss.n354 iovss.n353 0.818682
R650 iovss.n177 iovss.n176 0.818682
R651 iovss.n342 iovss.n341 0.818682
R652 iovss.n340 iovss.n184 0.818682
R653 iovss.n339 iovss.n338 0.818682
R654 iovss.n186 iovss.n185 0.818682
R655 iovss.n327 iovss.n326 0.818682
R656 iovss.n325 iovss.n193 0.818682
R657 iovss.n324 iovss.n323 0.818682
R658 iovss.n195 iovss.n194 0.818682
R659 iovss.n312 iovss.n311 0.818682
R660 iovss.n310 iovss.n202 0.818682
R661 iovss.n309 iovss.n308 0.818682
R662 iovss.n204 iovss.n203 0.818682
R663 iovss.n297 iovss.n296 0.818682
R664 iovss.n295 iovss.n211 0.818682
R665 iovss.n294 iovss.n293 0.818682
R666 iovss.n213 iovss.n212 0.818682
R667 iovss.n282 iovss.n281 0.818682
R668 iovss.n280 iovss.n220 0.818682
R669 iovss.n279 iovss.n278 0.818682
R670 iovss.n222 iovss.n221 0.818682
R671 iovss.n267 iovss.n266 0.818682
R672 iovss.n265 iovss.n229 0.818682
R673 iovss.n264 iovss.n263 0.818682
R674 iovss.n231 iovss.n230 0.818682
R675 iovss.n252 iovss.n251 0.818682
R676 iovss.n250 iovss.n238 0.818682
R677 iovss.n249 iovss.n248 0.818682
R678 iovss.n679 iovss.n98 0.818682
R679 iovss.n667 iovss.n666 0.818682
R680 iovss.n665 iovss.n476 0.818682
R681 iovss.n664 iovss.n663 0.818682
R682 iovss.n478 iovss.n477 0.818682
R683 iovss.n652 iovss.n651 0.818682
R684 iovss.n650 iovss.n485 0.818682
R685 iovss.n649 iovss.n648 0.818682
R686 iovss.n487 iovss.n486 0.818682
R687 iovss.n637 iovss.n636 0.818682
R688 iovss.n635 iovss.n494 0.818682
R689 iovss.n634 iovss.n633 0.818682
R690 iovss.n496 iovss.n495 0.818682
R691 iovss.n622 iovss.n621 0.818682
R692 iovss.n620 iovss.n503 0.818682
R693 iovss.n619 iovss.n618 0.818682
R694 iovss.n505 iovss.n504 0.818682
R695 iovss.n607 iovss.n606 0.818682
R696 iovss.n605 iovss.n512 0.818682
R697 iovss.n604 iovss.n603 0.818682
R698 iovss.n514 iovss.n513 0.818682
R699 iovss.n592 iovss.n591 0.818682
R700 iovss.n590 iovss.n521 0.818682
R701 iovss.n589 iovss.n588 0.818682
R702 iovss.n523 iovss.n522 0.818682
R703 iovss.n577 iovss.n576 0.818682
R704 iovss.n575 iovss.n530 0.818682
R705 iovss.n574 iovss.n573 0.818682
R706 iovss.n532 iovss.n531 0.818682
R707 iovss.n562 iovss.n561 0.818682
R708 iovss.n560 iovss.n539 0.818682
R709 iovss.n559 iovss.n558 0.818682
R710 iovss.n541 iovss.n540 0.818682
R711 iovss.n468 iovss.n72 0.818682
R712 iovss.n688 iovss.n687 0.818682
R713 iovss.n469 iovss.n458 0.818682
R714 iovss.n680 iovss.n113 0.818682
R715 iovss.n548 iovss.n547 0.818682
R716 iovss.n549 iovss.n541 0.818682
R717 iovss.n558 iovss.n557 0.818682
R718 iovss.n543 iovss.n539 0.818682
R719 iovss.n563 iovss.n562 0.818682
R720 iovss.n564 iovss.n532 0.818682
R721 iovss.n573 iovss.n572 0.818682
R722 iovss.n534 iovss.n530 0.818682
R723 iovss.n578 iovss.n577 0.818682
R724 iovss.n579 iovss.n523 0.818682
R725 iovss.n588 iovss.n587 0.818682
R726 iovss.n525 iovss.n521 0.818682
R727 iovss.n593 iovss.n592 0.818682
R728 iovss.n594 iovss.n514 0.818682
R729 iovss.n603 iovss.n602 0.818682
R730 iovss.n516 iovss.n512 0.818682
R731 iovss.n608 iovss.n607 0.818682
R732 iovss.n609 iovss.n505 0.818682
R733 iovss.n618 iovss.n617 0.818682
R734 iovss.n507 iovss.n503 0.818682
R735 iovss.n623 iovss.n622 0.818682
R736 iovss.n624 iovss.n496 0.818682
R737 iovss.n633 iovss.n632 0.818682
R738 iovss.n498 iovss.n494 0.818682
R739 iovss.n638 iovss.n637 0.818682
R740 iovss.n639 iovss.n487 0.818682
R741 iovss.n648 iovss.n647 0.818682
R742 iovss.n489 iovss.n485 0.818682
R743 iovss.n653 iovss.n652 0.818682
R744 iovss.n654 iovss.n478 0.818682
R745 iovss.n663 iovss.n662 0.818682
R746 iovss.n480 iovss.n476 0.818682
R747 iovss.n668 iovss.n667 0.818682
R748 iovss.n669 iovss.n468 0.818682
R749 iovss.n687 iovss.n686 0.818682
R750 iovss.n471 iovss.n469 0.818682
R751 iovss.n681 iovss.n680 0.818682
R752 iovss.n249 iovss.n239 0.416993
R753 iovss.n546 iovss.n540 0.416993
R754 iovss.n696 iovss 0.341436
R755 iovss.n243 iovss.n242 0.201704
R756 iovss.n552 iovss.n545 0.201704
R757 iovss.n883 iovss.n882 0.2005
R758 iovss.n167 iovss.n163 0.2005
R759 iovss.n878 iovss.n877 0.2005
R760 iovss.n366 iovss.n165 0.2005
R761 iovss.n365 iovss.n364 0.2005
R762 iovss.n174 iovss.n170 0.2005
R763 iovss.n360 iovss.n359 0.2005
R764 iovss.n351 iovss.n172 0.2005
R765 iovss.n350 iovss.n349 0.2005
R766 iovss.n183 iovss.n179 0.2005
R767 iovss.n345 iovss.n344 0.2005
R768 iovss.n336 iovss.n181 0.2005
R769 iovss.n335 iovss.n334 0.2005
R770 iovss.n192 iovss.n188 0.2005
R771 iovss.n330 iovss.n329 0.2005
R772 iovss.n321 iovss.n190 0.2005
R773 iovss.n320 iovss.n319 0.2005
R774 iovss.n201 iovss.n197 0.2005
R775 iovss.n315 iovss.n314 0.2005
R776 iovss.n306 iovss.n199 0.2005
R777 iovss.n305 iovss.n304 0.2005
R778 iovss.n210 iovss.n206 0.2005
R779 iovss.n300 iovss.n299 0.2005
R780 iovss.n291 iovss.n208 0.2005
R781 iovss.n290 iovss.n289 0.2005
R782 iovss.n219 iovss.n215 0.2005
R783 iovss.n285 iovss.n284 0.2005
R784 iovss.n276 iovss.n217 0.2005
R785 iovss.n275 iovss.n274 0.2005
R786 iovss.n228 iovss.n224 0.2005
R787 iovss.n270 iovss.n269 0.2005
R788 iovss.n261 iovss.n226 0.2005
R789 iovss.n260 iovss.n259 0.2005
R790 iovss.n237 iovss.n233 0.2005
R791 iovss.n255 iovss.n254 0.2005
R792 iovss.n246 iovss.n235 0.2005
R793 iovss.n245 iovss.n244 0.2005
R794 iovss.n678 iovss.n677 0.2005
R795 iovss.n683 iovss.n682 0.2005
R796 iovss.n685 iovss.n684 0.2005
R797 iovss.n472 iovss.n470 0.2005
R798 iovss.n671 iovss.n670 0.2005
R799 iovss.n475 iovss.n474 0.2005
R800 iovss.n661 iovss.n660 0.2005
R801 iovss.n481 iovss.n479 0.2005
R802 iovss.n656 iovss.n655 0.2005
R803 iovss.n484 iovss.n483 0.2005
R804 iovss.n646 iovss.n645 0.2005
R805 iovss.n490 iovss.n488 0.2005
R806 iovss.n641 iovss.n640 0.2005
R807 iovss.n493 iovss.n492 0.2005
R808 iovss.n631 iovss.n630 0.2005
R809 iovss.n499 iovss.n497 0.2005
R810 iovss.n626 iovss.n625 0.2005
R811 iovss.n502 iovss.n501 0.2005
R812 iovss.n616 iovss.n615 0.2005
R813 iovss.n508 iovss.n506 0.2005
R814 iovss.n611 iovss.n610 0.2005
R815 iovss.n511 iovss.n510 0.2005
R816 iovss.n601 iovss.n600 0.2005
R817 iovss.n517 iovss.n515 0.2005
R818 iovss.n596 iovss.n595 0.2005
R819 iovss.n520 iovss.n519 0.2005
R820 iovss.n586 iovss.n585 0.2005
R821 iovss.n526 iovss.n524 0.2005
R822 iovss.n581 iovss.n580 0.2005
R823 iovss.n529 iovss.n528 0.2005
R824 iovss.n571 iovss.n570 0.2005
R825 iovss.n535 iovss.n533 0.2005
R826 iovss.n566 iovss.n565 0.2005
R827 iovss.n538 iovss.n537 0.2005
R828 iovss.n556 iovss.n555 0.2005
R829 iovss.n544 iovss.n542 0.2005
R830 iovss.n551 iovss.n550 0.2005
R831 iovss.n778 iovss 0.1105
R832 iovss.n1016 iovss 0.1105
R833 iovss.n445 iovss 0.1105
R834 iovss.n882 iovss.n881 0.1105
R835 iovss.n880 iovss.n163 0.1105
R836 iovss.n879 iovss.n878 0.1105
R837 iovss.n165 iovss.n164 0.1105
R838 iovss.n364 iovss.n363 0.1105
R839 iovss.n362 iovss.n170 0.1105
R840 iovss.n361 iovss.n360 0.1105
R841 iovss.n172 iovss.n171 0.1105
R842 iovss.n349 iovss.n348 0.1105
R843 iovss.n347 iovss.n179 0.1105
R844 iovss.n346 iovss.n345 0.1105
R845 iovss.n181 iovss.n180 0.1105
R846 iovss.n334 iovss.n333 0.1105
R847 iovss.n332 iovss.n188 0.1105
R848 iovss.n331 iovss.n330 0.1105
R849 iovss.n190 iovss.n189 0.1105
R850 iovss.n319 iovss.n318 0.1105
R851 iovss.n317 iovss.n197 0.1105
R852 iovss.n316 iovss.n315 0.1105
R853 iovss.n199 iovss.n198 0.1105
R854 iovss.n304 iovss.n303 0.1105
R855 iovss.n302 iovss.n206 0.1105
R856 iovss.n301 iovss.n300 0.1105
R857 iovss.n208 iovss.n207 0.1105
R858 iovss.n289 iovss.n288 0.1105
R859 iovss.n287 iovss.n215 0.1105
R860 iovss.n286 iovss.n285 0.1105
R861 iovss.n217 iovss.n216 0.1105
R862 iovss.n274 iovss.n273 0.1105
R863 iovss.n272 iovss.n224 0.1105
R864 iovss.n271 iovss.n270 0.1105
R865 iovss.n226 iovss.n225 0.1105
R866 iovss.n259 iovss.n258 0.1105
R867 iovss.n257 iovss.n233 0.1105
R868 iovss.n256 iovss.n255 0.1105
R869 iovss.n235 iovss.n234 0.1105
R870 iovss.n677 iovss.n676 0.1105
R871 iovss.n683 iovss.n675 0.1105
R872 iovss.n684 iovss.n674 0.1105
R873 iovss.n673 iovss.n472 0.1105
R874 iovss.n672 iovss.n671 0.1105
R875 iovss.n474 iovss.n473 0.1105
R876 iovss.n660 iovss.n659 0.1105
R877 iovss.n658 iovss.n481 0.1105
R878 iovss.n657 iovss.n656 0.1105
R879 iovss.n483 iovss.n482 0.1105
R880 iovss.n645 iovss.n644 0.1105
R881 iovss.n643 iovss.n490 0.1105
R882 iovss.n642 iovss.n641 0.1105
R883 iovss.n492 iovss.n491 0.1105
R884 iovss.n630 iovss.n629 0.1105
R885 iovss.n628 iovss.n499 0.1105
R886 iovss.n627 iovss.n626 0.1105
R887 iovss.n501 iovss.n500 0.1105
R888 iovss.n615 iovss.n614 0.1105
R889 iovss.n613 iovss.n508 0.1105
R890 iovss.n612 iovss.n611 0.1105
R891 iovss.n510 iovss.n509 0.1105
R892 iovss.n600 iovss.n599 0.1105
R893 iovss.n598 iovss.n517 0.1105
R894 iovss.n597 iovss.n596 0.1105
R895 iovss.n519 iovss.n518 0.1105
R896 iovss.n585 iovss.n584 0.1105
R897 iovss.n583 iovss.n526 0.1105
R898 iovss.n582 iovss.n581 0.1105
R899 iovss.n528 iovss.n527 0.1105
R900 iovss.n570 iovss.n569 0.1105
R901 iovss.n568 iovss.n535 0.1105
R902 iovss.n567 iovss.n566 0.1105
R903 iovss.n537 iovss.n536 0.1105
R904 iovss.n555 iovss.n554 0.1105
R905 iovss.n553 iovss.n544 0.1105
R906 iovss.n553 iovss.n552 0.0568704
R907 iovss.n243 iovss.n234 0.0568704
R908 iovss.n120 iovss.n119 0.0432778
R909 iovss.n121 iovss.n120 0.0432778
R910 iovss.n122 iovss.n121 0.0432778
R911 iovss.n123 iovss.n122 0.0432778
R912 iovss.n124 iovss.n123 0.0432778
R913 iovss.n125 iovss.n124 0.0432778
R914 iovss.n897 iovss.n125 0.0432778
R915 iovss.n897 iovss.n896 0.0432778
R916 iovss.n896 iovss.n126 0.0432778
R917 iovss.n129 iovss.n126 0.0432778
R918 iovss.n130 iovss.n129 0.0432778
R919 iovss.n131 iovss.n130 0.0432778
R920 iovss.n132 iovss.n131 0.0432778
R921 iovss.n772 iovss.n132 0.0432778
R922 iovss.n773 iovss.n772 0.0432778
R923 iovss.n869 iovss.n773 0.0432778
R924 iovss.n869 iovss.n868 0.0432778
R925 iovss.n868 iovss.n866 0.0432778
R926 iovss.n866 iovss.n864 0.0432778
R927 iovss.n864 iovss.n862 0.0432778
R928 iovss.n862 iovss.n860 0.0432778
R929 iovss.n860 iovss.n858 0.0432778
R930 iovss.n858 iovss.n856 0.0432778
R931 iovss.n856 iovss.n854 0.0432778
R932 iovss.n854 iovss.n852 0.0432778
R933 iovss.n852 iovss.n850 0.0432778
R934 iovss.n850 iovss.n848 0.0432778
R935 iovss.n848 iovss.n846 0.0432778
R936 iovss.n846 iovss.n844 0.0432778
R937 iovss.n844 iovss.n842 0.0432778
R938 iovss.n842 iovss.n840 0.0432778
R939 iovss.n840 iovss.n838 0.0432778
R940 iovss.n838 iovss.n836 0.0432778
R941 iovss.n836 iovss.n834 0.0432778
R942 iovss.n834 iovss.n832 0.0432778
R943 iovss.n832 iovss.n830 0.0432778
R944 iovss.n830 iovss.n828 0.0432778
R945 iovss.n828 iovss.n826 0.0432778
R946 iovss.n826 iovss.n824 0.0432778
R947 iovss.n824 iovss.n822 0.0432778
R948 iovss.n822 iovss.n820 0.0432778
R949 iovss.n820 iovss.n818 0.0432778
R950 iovss.n818 iovss.n816 0.0432778
R951 iovss.n816 iovss.n814 0.0432778
R952 iovss.n814 iovss.n812 0.0432778
R953 iovss.n812 iovss.n810 0.0432778
R954 iovss.n810 iovss.n808 0.0432778
R955 iovss.n808 iovss.n806 0.0432778
R956 iovss.n806 iovss.n804 0.0432778
R957 iovss.n804 iovss.n802 0.0432778
R958 iovss.n802 iovss.n800 0.0432778
R959 iovss.n800 iovss.n798 0.0432778
R960 iovss.n798 iovss.n796 0.0432778
R961 iovss.n796 iovss.n794 0.0432778
R962 iovss.n794 iovss.n792 0.0432778
R963 iovss.n792 iovss.n790 0.0432778
R964 iovss.n790 iovss.n788 0.0432778
R965 iovss.n788 iovss.n786 0.0432778
R966 iovss.n786 iovss.n784 0.0432778
R967 iovss.n784 iovss.n782 0.0432778
R968 iovss.n782 iovss.n780 0.0432778
R969 iovss.n89 iovss.n83 0.0432778
R970 iovss.n89 iovss.n88 0.0432778
R971 iovss.n88 iovss.n87 0.0432778
R972 iovss.n87 iovss.n86 0.0432778
R973 iovss.n86 iovss.n85 0.0432778
R974 iovss.n85 iovss.n84 0.0432778
R975 iovss.n84 iovss.n63 0.0432778
R976 iovss.n908 iovss.n63 0.0432778
R977 iovss.n909 iovss.n908 0.0432778
R978 iovss.n910 iovss.n909 0.0432778
R979 iovss.n910 iovss.n59 0.0432778
R980 iovss.n917 iovss.n59 0.0432778
R981 iovss.n918 iovss.n917 0.0432778
R982 iovss.n999 iovss.n918 0.0432778
R983 iovss.n999 iovss.n998 0.0432778
R984 iovss.n998 iovss.n996 0.0432778
R985 iovss.n996 iovss.n994 0.0432778
R986 iovss.n994 iovss.n992 0.0432778
R987 iovss.n992 iovss.n990 0.0432778
R988 iovss.n990 iovss.n988 0.0432778
R989 iovss.n988 iovss.n986 0.0432778
R990 iovss.n986 iovss.n984 0.0432778
R991 iovss.n984 iovss.n982 0.0432778
R992 iovss.n982 iovss.n980 0.0432778
R993 iovss.n980 iovss.n978 0.0432778
R994 iovss.n978 iovss.n976 0.0432778
R995 iovss.n976 iovss.n974 0.0432778
R996 iovss.n974 iovss.n972 0.0432778
R997 iovss.n972 iovss.n970 0.0432778
R998 iovss.n970 iovss.n968 0.0432778
R999 iovss.n968 iovss.n966 0.0432778
R1000 iovss.n966 iovss.n964 0.0432778
R1001 iovss.n964 iovss.n962 0.0432778
R1002 iovss.n962 iovss.n960 0.0432778
R1003 iovss.n960 iovss.n958 0.0432778
R1004 iovss.n958 iovss.n956 0.0432778
R1005 iovss.n956 iovss.n954 0.0432778
R1006 iovss.n954 iovss.n952 0.0432778
R1007 iovss.n952 iovss.n950 0.0432778
R1008 iovss.n950 iovss.n948 0.0432778
R1009 iovss.n948 iovss.n946 0.0432778
R1010 iovss.n946 iovss.n944 0.0432778
R1011 iovss.n944 iovss.n942 0.0432778
R1012 iovss.n942 iovss.n940 0.0432778
R1013 iovss.n940 iovss.n938 0.0432778
R1014 iovss.n938 iovss.n936 0.0432778
R1015 iovss.n936 iovss.n934 0.0432778
R1016 iovss.n934 iovss.n932 0.0432778
R1017 iovss.n932 iovss.n930 0.0432778
R1018 iovss.n930 iovss.n928 0.0432778
R1019 iovss.n928 iovss.n926 0.0432778
R1020 iovss.n926 iovss.n924 0.0432778
R1021 iovss.n924 iovss.n922 0.0432778
R1022 iovss.n922 iovss.n920 0.0432778
R1023 iovss.n920 iovss.n35 0.0432778
R1024 iovss.n1004 iovss.n35 0.0432778
R1025 iovss.n1006 iovss.n1004 0.0432778
R1026 iovss.n1007 iovss.n1006 0.0432778
R1027 iovss.n1007 iovss.n8 0.0432778
R1028 iovss.n1014 iovss.n8 0.0432778
R1029 iovss.n1015 iovss.n1014 0.0432778
R1030 iovss.n893 iovss.n892 0.0347222
R1031 iovss.n892 iovss.n891 0.0347222
R1032 iovss.n891 iovss.n128 0.0347222
R1033 iovss.n887 iovss.n128 0.0347222
R1034 iovss.n704 iovss.n703 0.0347222
R1035 iovss.n705 iovss.n704 0.0347222
R1036 iovss.n705 iovss.n446 0.0347222
R1037 iovss.n711 iovss.n446 0.0347222
R1038 iovss.n912 iovss.n61 0.0347222
R1039 iovss.n913 iovss.n912 0.0347222
R1040 iovss.n915 iovss.n913 0.0347222
R1041 iovss.n915 iovss.n914 0.0347222
R1042 iovss.n907 iovss.n62 0.0347222
R1043 iovss.n911 iovss.n62 0.0347222
R1044 iovss.n911 iovss.n60 0.0347222
R1045 iovss.n916 iovss.n60 0.0347222
R1046 iovss.n916 iovss.n58 0.0347222
R1047 iovss.n1000 iovss.n58 0.0347222
R1048 iovss.n1013 iovss.n4 0.0347222
R1049 iovss.n1017 iovss.n4 0.0347222
R1050 iovss.n702 iovss.n700 0.0347222
R1051 iovss.n706 iovss.n447 0.0347222
R1052 iovss.n710 iovss.n708 0.0347222
R1053 iovss.n895 iovss.n894 0.0347222
R1054 iovss.n894 iovss.n127 0.0347222
R1055 iovss.n890 iovss.n127 0.0347222
R1056 iovss.n890 iovss.n889 0.0347222
R1057 iovss.n889 iovss.n888 0.0347222
R1058 iovss.n888 iovss.n133 0.0347222
R1059 iovss.n119 iovss.n1 0.0231984
R1060 iovss.n83 iovss.n1 0.0231984
R1061 iovss.n112 iovss.n1 0.0205794
R1062 iovss.n695 iovss.n1 0.0205794
R1063 iovss.n94 iovss.n67 0.0180786
R1064 iovss.n93 iovss.n91 0.0180786
R1065 iovss.n92 iovss.n68 0.0180786
R1066 iovss.n90 iovss.n81 0.0180786
R1067 iovss.n82 iovss.n69 0.0180786
R1068 iovss.n80 iovss.n78 0.0180786
R1069 iovss.n79 iovss.n70 0.0180786
R1070 iovss.n77 iovss.n75 0.0180786
R1071 iovss.n76 iovss.n71 0.0180786
R1072 iovss.n74 iovss.n73 0.0180786
R1073 iovss.n907 iovss.n64 0.0180786
R1074 iovss.n1000 iovss.n12 0.0180786
R1075 iovss.n997 iovss.n37 0.0180786
R1076 iovss.n995 iovss.n13 0.0180786
R1077 iovss.n993 iovss.n38 0.0180786
R1078 iovss.n991 iovss.n14 0.0180786
R1079 iovss.n989 iovss.n39 0.0180786
R1080 iovss.n987 iovss.n15 0.0180786
R1081 iovss.n985 iovss.n40 0.0180786
R1082 iovss.n983 iovss.n16 0.0180786
R1083 iovss.n981 iovss.n41 0.0180786
R1084 iovss.n979 iovss.n17 0.0180786
R1085 iovss.n977 iovss.n42 0.0180786
R1086 iovss.n975 iovss.n18 0.0180786
R1087 iovss.n973 iovss.n43 0.0180786
R1088 iovss.n971 iovss.n19 0.0180786
R1089 iovss.n969 iovss.n44 0.0180786
R1090 iovss.n967 iovss.n20 0.0180786
R1091 iovss.n965 iovss.n45 0.0180786
R1092 iovss.n963 iovss.n21 0.0180786
R1093 iovss.n961 iovss.n46 0.0180786
R1094 iovss.n959 iovss.n22 0.0180786
R1095 iovss.n957 iovss.n47 0.0180786
R1096 iovss.n955 iovss.n23 0.0180786
R1097 iovss.n953 iovss.n48 0.0180786
R1098 iovss.n951 iovss.n24 0.0180786
R1099 iovss.n949 iovss.n49 0.0180786
R1100 iovss.n947 iovss.n25 0.0180786
R1101 iovss.n945 iovss.n50 0.0180786
R1102 iovss.n943 iovss.n26 0.0180786
R1103 iovss.n941 iovss.n51 0.0180786
R1104 iovss.n939 iovss.n27 0.0180786
R1105 iovss.n937 iovss.n52 0.0180786
R1106 iovss.n935 iovss.n28 0.0180786
R1107 iovss.n933 iovss.n53 0.0180786
R1108 iovss.n931 iovss.n29 0.0180786
R1109 iovss.n929 iovss.n54 0.0180786
R1110 iovss.n927 iovss.n30 0.0180786
R1111 iovss.n925 iovss.n55 0.0180786
R1112 iovss.n923 iovss.n31 0.0180786
R1113 iovss.n921 iovss.n56 0.0180786
R1114 iovss.n919 iovss.n32 0.0180786
R1115 iovss.n1002 iovss.n36 0.0180786
R1116 iovss.n1003 iovss.n33 0.0180786
R1117 iovss.n1005 iovss.n34 0.0180786
R1118 iovss.n1010 iovss.n1008 0.0180786
R1119 iovss.n1009 iovss.n9 0.0180786
R1120 iovss.n1017 iovss.n7 0.0180786
R1121 iovss.n1013 iovss.n9 0.0180786
R1122 iovss.n1010 iovss.n1009 0.0180786
R1123 iovss.n1008 iovss.n34 0.0180786
R1124 iovss.n1005 iovss.n33 0.0180786
R1125 iovss.n1003 iovss.n1002 0.0180786
R1126 iovss.n36 iovss.n32 0.0180786
R1127 iovss.n919 iovss.n56 0.0180786
R1128 iovss.n921 iovss.n31 0.0180786
R1129 iovss.n923 iovss.n55 0.0180786
R1130 iovss.n925 iovss.n30 0.0180786
R1131 iovss.n927 iovss.n54 0.0180786
R1132 iovss.n929 iovss.n29 0.0180786
R1133 iovss.n931 iovss.n53 0.0180786
R1134 iovss.n933 iovss.n28 0.0180786
R1135 iovss.n935 iovss.n52 0.0180786
R1136 iovss.n937 iovss.n27 0.0180786
R1137 iovss.n939 iovss.n51 0.0180786
R1138 iovss.n941 iovss.n26 0.0180786
R1139 iovss.n943 iovss.n50 0.0180786
R1140 iovss.n945 iovss.n25 0.0180786
R1141 iovss.n947 iovss.n49 0.0180786
R1142 iovss.n949 iovss.n24 0.0180786
R1143 iovss.n951 iovss.n48 0.0180786
R1144 iovss.n953 iovss.n23 0.0180786
R1145 iovss.n955 iovss.n47 0.0180786
R1146 iovss.n957 iovss.n22 0.0180786
R1147 iovss.n959 iovss.n46 0.0180786
R1148 iovss.n961 iovss.n21 0.0180786
R1149 iovss.n963 iovss.n45 0.0180786
R1150 iovss.n965 iovss.n20 0.0180786
R1151 iovss.n967 iovss.n44 0.0180786
R1152 iovss.n969 iovss.n19 0.0180786
R1153 iovss.n971 iovss.n43 0.0180786
R1154 iovss.n973 iovss.n18 0.0180786
R1155 iovss.n975 iovss.n42 0.0180786
R1156 iovss.n977 iovss.n17 0.0180786
R1157 iovss.n979 iovss.n41 0.0180786
R1158 iovss.n981 iovss.n16 0.0180786
R1159 iovss.n983 iovss.n40 0.0180786
R1160 iovss.n985 iovss.n15 0.0180786
R1161 iovss.n987 iovss.n39 0.0180786
R1162 iovss.n989 iovss.n14 0.0180786
R1163 iovss.n991 iovss.n38 0.0180786
R1164 iovss.n993 iovss.n13 0.0180786
R1165 iovss.n995 iovss.n37 0.0180786
R1166 iovss.n997 iovss.n12 0.0180786
R1167 iovss.n7 iovss.n3 0.0180786
R1168 iovss.n453 iovss.n451 0.0180786
R1169 iovss.n698 iovss.n693 0.0180786
R1170 iovss.n694 iovss.n454 0.0180786
R1171 iovss.n466 iovss.n455 0.0180786
R1172 iovss.n691 iovss.n456 0.0180786
R1173 iovss.n463 iovss.n461 0.0180786
R1174 iovss.n460 iovss.n459 0.0180786
R1175 iovss.n712 iovss.n371 0.0180786
R1176 iovss.n713 iovss.n372 0.0180786
R1177 iovss.n714 iovss.n373 0.0180786
R1178 iovss.n715 iovss.n374 0.0180786
R1179 iovss.n716 iovss.n375 0.0180786
R1180 iovss.n717 iovss.n376 0.0180786
R1181 iovss.n718 iovss.n377 0.0180786
R1182 iovss.n719 iovss.n378 0.0180786
R1183 iovss.n720 iovss.n379 0.0180786
R1184 iovss.n721 iovss.n380 0.0180786
R1185 iovss.n722 iovss.n381 0.0180786
R1186 iovss.n723 iovss.n382 0.0180786
R1187 iovss.n724 iovss.n383 0.0180786
R1188 iovss.n725 iovss.n384 0.0180786
R1189 iovss.n726 iovss.n385 0.0180786
R1190 iovss.n727 iovss.n386 0.0180786
R1191 iovss.n728 iovss.n387 0.0180786
R1192 iovss.n729 iovss.n388 0.0180786
R1193 iovss.n730 iovss.n389 0.0180786
R1194 iovss.n731 iovss.n390 0.0180786
R1195 iovss.n732 iovss.n391 0.0180786
R1196 iovss.n733 iovss.n392 0.0180786
R1197 iovss.n734 iovss.n393 0.0180786
R1198 iovss.n735 iovss.n394 0.0180786
R1199 iovss.n743 iovss.n394 0.0180786
R1200 iovss.n746 iovss.n443 0.0180786
R1201 iovss.n735 iovss.n396 0.0180786
R1202 iovss.n734 iovss.n398 0.0180786
R1203 iovss.n733 iovss.n400 0.0180786
R1204 iovss.n732 iovss.n402 0.0180786
R1205 iovss.n731 iovss.n404 0.0180786
R1206 iovss.n730 iovss.n406 0.0180786
R1207 iovss.n729 iovss.n408 0.0180786
R1208 iovss.n728 iovss.n410 0.0180786
R1209 iovss.n727 iovss.n412 0.0180786
R1210 iovss.n726 iovss.n414 0.0180786
R1211 iovss.n725 iovss.n416 0.0180786
R1212 iovss.n724 iovss.n418 0.0180786
R1213 iovss.n723 iovss.n420 0.0180786
R1214 iovss.n722 iovss.n422 0.0180786
R1215 iovss.n721 iovss.n424 0.0180786
R1216 iovss.n720 iovss.n426 0.0180786
R1217 iovss.n719 iovss.n428 0.0180786
R1218 iovss.n718 iovss.n430 0.0180786
R1219 iovss.n717 iovss.n432 0.0180786
R1220 iovss.n716 iovss.n434 0.0180786
R1221 iovss.n715 iovss.n436 0.0180786
R1222 iovss.n714 iovss.n438 0.0180786
R1223 iovss.n713 iovss.n440 0.0180786
R1224 iovss.n712 iovss.n441 0.0180786
R1225 iovss.n744 iovss.n743 0.0180786
R1226 iovss.n744 iovss.n443 0.0180786
R1227 iovss.n99 iovss.n97 0.0180786
R1228 iovss.n901 iovss.n111 0.0180786
R1229 iovss.n900 iovss.n100 0.0180786
R1230 iovss.n110 iovss.n109 0.0180786
R1231 iovss.n114 iovss.n101 0.0180786
R1232 iovss.n108 iovss.n107 0.0180786
R1233 iovss.n115 iovss.n102 0.0180786
R1234 iovss.n106 iovss.n105 0.0180786
R1235 iovss.n116 iovss.n103 0.0180786
R1236 iovss.n898 iovss.n118 0.0180786
R1237 iovss.n895 iovss.n104 0.0180786
R1238 iovss.n771 iovss.n136 0.0180786
R1239 iovss.n871 iovss.n870 0.0180786
R1240 iovss.n867 iovss.n137 0.0180786
R1241 iovss.n865 iovss.n770 0.0180786
R1242 iovss.n863 iovss.n138 0.0180786
R1243 iovss.n861 iovss.n769 0.0180786
R1244 iovss.n859 iovss.n139 0.0180786
R1245 iovss.n857 iovss.n768 0.0180786
R1246 iovss.n855 iovss.n140 0.0180786
R1247 iovss.n853 iovss.n767 0.0180786
R1248 iovss.n851 iovss.n141 0.0180786
R1249 iovss.n849 iovss.n766 0.0180786
R1250 iovss.n847 iovss.n142 0.0180786
R1251 iovss.n845 iovss.n765 0.0180786
R1252 iovss.n843 iovss.n143 0.0180786
R1253 iovss.n841 iovss.n764 0.0180786
R1254 iovss.n839 iovss.n144 0.0180786
R1255 iovss.n837 iovss.n763 0.0180786
R1256 iovss.n835 iovss.n145 0.0180786
R1257 iovss.n833 iovss.n762 0.0180786
R1258 iovss.n831 iovss.n146 0.0180786
R1259 iovss.n829 iovss.n761 0.0180786
R1260 iovss.n827 iovss.n147 0.0180786
R1261 iovss.n825 iovss.n760 0.0180786
R1262 iovss.n823 iovss.n148 0.0180786
R1263 iovss.n821 iovss.n759 0.0180786
R1264 iovss.n819 iovss.n149 0.0180786
R1265 iovss.n817 iovss.n758 0.0180786
R1266 iovss.n815 iovss.n150 0.0180786
R1267 iovss.n813 iovss.n757 0.0180786
R1268 iovss.n811 iovss.n151 0.0180786
R1269 iovss.n809 iovss.n756 0.0180786
R1270 iovss.n807 iovss.n152 0.0180786
R1271 iovss.n805 iovss.n755 0.0180786
R1272 iovss.n803 iovss.n153 0.0180786
R1273 iovss.n801 iovss.n754 0.0180786
R1274 iovss.n799 iovss.n154 0.0180786
R1275 iovss.n797 iovss.n753 0.0180786
R1276 iovss.n795 iovss.n155 0.0180786
R1277 iovss.n793 iovss.n752 0.0180786
R1278 iovss.n791 iovss.n156 0.0180786
R1279 iovss.n789 iovss.n751 0.0180786
R1280 iovss.n787 iovss.n157 0.0180786
R1281 iovss.n785 iovss.n750 0.0180786
R1282 iovss.n783 iovss.n158 0.0180786
R1283 iovss.n781 iovss.n749 0.0180786
R1284 iovss.n779 iovss.n159 0.0180786
R1285 iovss.n779 iovss.n748 0.0180786
R1286 iovss.n776 iovss.n135 0.0180786
R1287 iovss.n777 iovss.n776 0.0180786
R1288 iovss.n781 iovss.n159 0.0180786
R1289 iovss.n783 iovss.n749 0.0180786
R1290 iovss.n785 iovss.n158 0.0180786
R1291 iovss.n787 iovss.n750 0.0180786
R1292 iovss.n789 iovss.n157 0.0180786
R1293 iovss.n791 iovss.n751 0.0180786
R1294 iovss.n793 iovss.n156 0.0180786
R1295 iovss.n795 iovss.n752 0.0180786
R1296 iovss.n797 iovss.n155 0.0180786
R1297 iovss.n799 iovss.n753 0.0180786
R1298 iovss.n801 iovss.n154 0.0180786
R1299 iovss.n803 iovss.n754 0.0180786
R1300 iovss.n805 iovss.n153 0.0180786
R1301 iovss.n807 iovss.n755 0.0180786
R1302 iovss.n809 iovss.n152 0.0180786
R1303 iovss.n811 iovss.n756 0.0180786
R1304 iovss.n813 iovss.n151 0.0180786
R1305 iovss.n815 iovss.n757 0.0180786
R1306 iovss.n817 iovss.n150 0.0180786
R1307 iovss.n819 iovss.n758 0.0180786
R1308 iovss.n821 iovss.n149 0.0180786
R1309 iovss.n823 iovss.n759 0.0180786
R1310 iovss.n825 iovss.n148 0.0180786
R1311 iovss.n827 iovss.n760 0.0180786
R1312 iovss.n829 iovss.n147 0.0180786
R1313 iovss.n831 iovss.n761 0.0180786
R1314 iovss.n833 iovss.n146 0.0180786
R1315 iovss.n835 iovss.n762 0.0180786
R1316 iovss.n837 iovss.n145 0.0180786
R1317 iovss.n839 iovss.n763 0.0180786
R1318 iovss.n841 iovss.n144 0.0180786
R1319 iovss.n843 iovss.n764 0.0180786
R1320 iovss.n845 iovss.n143 0.0180786
R1321 iovss.n847 iovss.n765 0.0180786
R1322 iovss.n849 iovss.n142 0.0180786
R1323 iovss.n851 iovss.n766 0.0180786
R1324 iovss.n853 iovss.n141 0.0180786
R1325 iovss.n855 iovss.n767 0.0180786
R1326 iovss.n857 iovss.n140 0.0180786
R1327 iovss.n859 iovss.n768 0.0180786
R1328 iovss.n861 iovss.n139 0.0180786
R1329 iovss.n863 iovss.n769 0.0180786
R1330 iovss.n865 iovss.n138 0.0180786
R1331 iovss.n867 iovss.n770 0.0180786
R1332 iovss.n870 iovss.n137 0.0180786
R1333 iovss.n871 iovss.n771 0.0180786
R1334 iovss.n136 iovss.n133 0.0180786
R1335 iovss.n748 iovss.n135 0.0180786
R1336 iovss.n898 iovss.n104 0.0180786
R1337 iovss.n118 iovss.n103 0.0180786
R1338 iovss.n116 iovss.n106 0.0180786
R1339 iovss.n105 iovss.n102 0.0180786
R1340 iovss.n115 iovss.n108 0.0180786
R1341 iovss.n107 iovss.n101 0.0180786
R1342 iovss.n114 iovss.n110 0.0180786
R1343 iovss.n109 iovss.n100 0.0180786
R1344 iovss.n901 iovss.n900 0.0180786
R1345 iovss.n111 iovss.n99 0.0180786
R1346 iovss.n903 iovss.n97 0.0180786
R1347 iovss.n459 iovss.n457 0.0180786
R1348 iovss.n461 iovss.n456 0.0180786
R1349 iovss.n691 iovss.n690 0.0180786
R1350 iovss.n467 iovss.n466 0.0180786
R1351 iovss.n698 iovss.n694 0.0180786
R1352 iovss.n693 iovss.n453 0.0180786
R1353 iovss.n451 iovss.n95 0.0180786
R1354 iovss.n74 iovss.n64 0.0180786
R1355 iovss.n73 iovss.n71 0.0180786
R1356 iovss.n77 iovss.n76 0.0180786
R1357 iovss.n75 iovss.n70 0.0180786
R1358 iovss.n80 iovss.n79 0.0180786
R1359 iovss.n78 iovss.n69 0.0180786
R1360 iovss.n90 iovss.n82 0.0180786
R1361 iovss.n81 iovss.n68 0.0180786
R1362 iovss.n93 iovss.n92 0.0180786
R1363 iovss.n91 iovss.n67 0.0180786
R1364 iovss.n905 iovss.n94 0.0180786
R1365 iovss.n425 iovss.n378 0.0180349
R1366 iovss.n434 iovss.n433 0.0180327
R1367 iovss.n400 iovss.n399 0.0180327
R1368 iovss.n416 iovss.n415 0.0180322
R1369 iovss.n462 iovss.n457 0.0180322
R1370 iovss.n710 iovss.n709 0.0180306
R1371 iovss.n407 iovss.n387 0.0180306
R1372 iovss.n707 iovss.n706 0.0180294
R1373 iovss.n409 iovss.n386 0.0180294
R1374 iovss.n418 iovss.n417 0.0180284
R1375 iovss.n432 iovss.n431 0.0180266
R1376 iovss.n398 iovss.n397 0.0180266
R1377 iovss.n689 iovss.n455 0.0180266
R1378 iovss.n423 iovss.n379 0.0180262
R1379 iovss.n436 iovss.n435 0.0180241
R1380 iovss.n402 iovss.n401 0.0180241
R1381 iovss.n427 iovss.n377 0.0180239
R1382 iovss.n439 iovss.n371 0.0180219
R1383 iovss.n405 iovss.n388 0.0180219
R1384 iovss.n414 iovss.n413 0.0180211
R1385 iovss.n700 iovss.n449 0.0180211
R1386 iovss.n420 iovss.n419 0.0180197
R1387 iovss.n702 iovss.n701 0.0180184
R1388 iovss.n411 iovss.n385 0.0180184
R1389 iovss.n421 iovss.n380 0.0180175
R1390 iovss.n465 iovss.n454 0.0180156
R1391 iovss.n430 iovss.n429 0.0180156
R1392 iovss.n396 iovss.n395 0.0180156
R1393 iovss.n438 iovss.n437 0.0180153
R1394 iovss.n404 iovss.n403 0.0180153
R1395 iovss.n437 iovss.n372 0.0180132
R1396 iovss.n403 iovss.n389 0.0180132
R1397 iovss.n429 iovss.n376 0.0180129
R1398 iovss.n395 iovss.n393 0.0180129
R1399 iovss.n467 iovss.n465 0.0180129
R1400 iovss.n422 iovss.n421 0.018011
R1401 iovss.n701 iovss.n447 0.0180101
R1402 iovss.n412 iovss.n411 0.0180101
R1403 iovss.n419 iovss.n381 0.0180088
R1404 iovss.n413 iovss.n384 0.0180073
R1405 iovss.n460 iovss.n449 0.0180073
R1406 iovss.n440 iovss.n439 0.0180066
R1407 iovss.n406 iovss.n405 0.0180066
R1408 iovss.n428 iovss.n427 0.0180046
R1409 iovss.n435 iovss.n373 0.0180044
R1410 iovss.n401 iovss.n390 0.0180044
R1411 iovss.n424 iovss.n423 0.0180022
R1412 iovss.n431 iovss.n375 0.0180018
R1413 iovss.n397 iovss.n392 0.0180018
R1414 iovss.n690 iovss.n689 0.0180018
R1415 iovss.n417 iovss.n382 0.0180001
R1416 iovss.n708 iovss.n707 0.017999
R1417 iovss.n410 iovss.n409 0.017999
R1418 iovss.n709 iovss.n441 0.0179979
R1419 iovss.n408 iovss.n407 0.0179979
R1420 iovss.n415 iovss.n383 0.0179962
R1421 iovss.n463 iovss.n462 0.0179962
R1422 iovss.n433 iovss.n374 0.0179957
R1423 iovss.n399 iovss.n391 0.0179957
R1424 iovss.n426 iovss.n425 0.0179935
R1425 iovss.n775 iovss 0.0127222
R1426 iovss.n696 iovss.n112 0.00748413
R1427 iovss.n780 iovss.n778 0.00748413
R1428 iovss.n696 iovss.n695 0.00748413
R1429 iovss.n1016 iovss.n1015 0.00748413
R1430 iovss.n248 iovss.n240 0.00740196
R1431 iovss.n248 iovss.n238 0.00740196
R1432 iovss.n252 iovss.n238 0.00740196
R1433 iovss.n252 iovss.n231 0.00740196
R1434 iovss.n263 iovss.n231 0.00740196
R1435 iovss.n263 iovss.n229 0.00740196
R1436 iovss.n267 iovss.n229 0.00740196
R1437 iovss.n267 iovss.n222 0.00740196
R1438 iovss.n278 iovss.n222 0.00740196
R1439 iovss.n278 iovss.n220 0.00740196
R1440 iovss.n282 iovss.n220 0.00740196
R1441 iovss.n282 iovss.n213 0.00740196
R1442 iovss.n293 iovss.n213 0.00740196
R1443 iovss.n293 iovss.n211 0.00740196
R1444 iovss.n297 iovss.n211 0.00740196
R1445 iovss.n297 iovss.n204 0.00740196
R1446 iovss.n308 iovss.n204 0.00740196
R1447 iovss.n308 iovss.n202 0.00740196
R1448 iovss.n312 iovss.n202 0.00740196
R1449 iovss.n312 iovss.n195 0.00740196
R1450 iovss.n323 iovss.n195 0.00740196
R1451 iovss.n323 iovss.n193 0.00740196
R1452 iovss.n327 iovss.n193 0.00740196
R1453 iovss.n327 iovss.n186 0.00740196
R1454 iovss.n338 iovss.n186 0.00740196
R1455 iovss.n338 iovss.n184 0.00740196
R1456 iovss.n342 iovss.n184 0.00740196
R1457 iovss.n342 iovss.n177 0.00740196
R1458 iovss.n353 iovss.n177 0.00740196
R1459 iovss.n353 iovss.n175 0.00740196
R1460 iovss.n357 iovss.n175 0.00740196
R1461 iovss.n357 iovss.n168 0.00740196
R1462 iovss.n368 iovss.n168 0.00740196
R1463 iovss.n369 iovss.n368 0.00740196
R1464 iovss.n875 iovss.n369 0.00740196
R1465 iovss.n875 iovss.n161 0.00740196
R1466 iovss.n884 iovss.n161 0.00740196
R1467 iovss.n250 iovss.n249 0.00740196
R1468 iovss.n251 iovss.n250 0.00740196
R1469 iovss.n251 iovss.n230 0.00740196
R1470 iovss.n264 iovss.n230 0.00740196
R1471 iovss.n265 iovss.n264 0.00740196
R1472 iovss.n266 iovss.n265 0.00740196
R1473 iovss.n266 iovss.n221 0.00740196
R1474 iovss.n279 iovss.n221 0.00740196
R1475 iovss.n280 iovss.n279 0.00740196
R1476 iovss.n281 iovss.n280 0.00740196
R1477 iovss.n281 iovss.n212 0.00740196
R1478 iovss.n294 iovss.n212 0.00740196
R1479 iovss.n295 iovss.n294 0.00740196
R1480 iovss.n296 iovss.n295 0.00740196
R1481 iovss.n296 iovss.n203 0.00740196
R1482 iovss.n309 iovss.n203 0.00740196
R1483 iovss.n310 iovss.n309 0.00740196
R1484 iovss.n311 iovss.n310 0.00740196
R1485 iovss.n311 iovss.n194 0.00740196
R1486 iovss.n324 iovss.n194 0.00740196
R1487 iovss.n325 iovss.n324 0.00740196
R1488 iovss.n326 iovss.n325 0.00740196
R1489 iovss.n326 iovss.n185 0.00740196
R1490 iovss.n339 iovss.n185 0.00740196
R1491 iovss.n340 iovss.n339 0.00740196
R1492 iovss.n341 iovss.n340 0.00740196
R1493 iovss.n341 iovss.n176 0.00740196
R1494 iovss.n354 iovss.n176 0.00740196
R1495 iovss.n355 iovss.n354 0.00740196
R1496 iovss.n356 iovss.n355 0.00740196
R1497 iovss.n356 iovss.n11 0.00740196
R1498 iovss.n741 iovss.n57 0.00740196
R1499 iovss.n874 iovss.n873 0.00740196
R1500 iovss.n559 iovss.n540 0.00740196
R1501 iovss.n560 iovss.n559 0.00740196
R1502 iovss.n561 iovss.n560 0.00740196
R1503 iovss.n561 iovss.n531 0.00740196
R1504 iovss.n574 iovss.n531 0.00740196
R1505 iovss.n575 iovss.n574 0.00740196
R1506 iovss.n576 iovss.n575 0.00740196
R1507 iovss.n576 iovss.n522 0.00740196
R1508 iovss.n589 iovss.n522 0.00740196
R1509 iovss.n590 iovss.n589 0.00740196
R1510 iovss.n591 iovss.n590 0.00740196
R1511 iovss.n591 iovss.n513 0.00740196
R1512 iovss.n604 iovss.n513 0.00740196
R1513 iovss.n605 iovss.n604 0.00740196
R1514 iovss.n606 iovss.n605 0.00740196
R1515 iovss.n606 iovss.n504 0.00740196
R1516 iovss.n619 iovss.n504 0.00740196
R1517 iovss.n620 iovss.n619 0.00740196
R1518 iovss.n621 iovss.n620 0.00740196
R1519 iovss.n621 iovss.n495 0.00740196
R1520 iovss.n634 iovss.n495 0.00740196
R1521 iovss.n635 iovss.n634 0.00740196
R1522 iovss.n636 iovss.n635 0.00740196
R1523 iovss.n636 iovss.n486 0.00740196
R1524 iovss.n649 iovss.n486 0.00740196
R1525 iovss.n650 iovss.n649 0.00740196
R1526 iovss.n651 iovss.n650 0.00740196
R1527 iovss.n651 iovss.n477 0.00740196
R1528 iovss.n664 iovss.n477 0.00740196
R1529 iovss.n665 iovss.n664 0.00740196
R1530 iovss.n666 iovss.n665 0.00740196
R1531 iovss.n688 iovss.n72 0.00740196
R1532 iovss.n458 iovss.n113 0.00740196
R1533 iovss.n547 iovss.n541 0.00740196
R1534 iovss.n558 iovss.n541 0.00740196
R1535 iovss.n558 iovss.n539 0.00740196
R1536 iovss.n562 iovss.n539 0.00740196
R1537 iovss.n562 iovss.n532 0.00740196
R1538 iovss.n573 iovss.n532 0.00740196
R1539 iovss.n573 iovss.n530 0.00740196
R1540 iovss.n577 iovss.n530 0.00740196
R1541 iovss.n577 iovss.n523 0.00740196
R1542 iovss.n588 iovss.n523 0.00740196
R1543 iovss.n588 iovss.n521 0.00740196
R1544 iovss.n592 iovss.n521 0.00740196
R1545 iovss.n592 iovss.n514 0.00740196
R1546 iovss.n603 iovss.n514 0.00740196
R1547 iovss.n603 iovss.n512 0.00740196
R1548 iovss.n607 iovss.n512 0.00740196
R1549 iovss.n607 iovss.n505 0.00740196
R1550 iovss.n618 iovss.n505 0.00740196
R1551 iovss.n618 iovss.n503 0.00740196
R1552 iovss.n622 iovss.n503 0.00740196
R1553 iovss.n622 iovss.n496 0.00740196
R1554 iovss.n633 iovss.n496 0.00740196
R1555 iovss.n633 iovss.n494 0.00740196
R1556 iovss.n637 iovss.n494 0.00740196
R1557 iovss.n637 iovss.n487 0.00740196
R1558 iovss.n648 iovss.n487 0.00740196
R1559 iovss.n648 iovss.n485 0.00740196
R1560 iovss.n652 iovss.n485 0.00740196
R1561 iovss.n652 iovss.n478 0.00740196
R1562 iovss.n663 iovss.n478 0.00740196
R1563 iovss.n663 iovss.n476 0.00740196
R1564 iovss.n667 iovss.n476 0.00740196
R1565 iovss.n667 iovss.n468 0.00740196
R1566 iovss.n687 iovss.n468 0.00740196
R1567 iovss.n687 iovss.n469 0.00740196
R1568 iovss.n680 iovss.n469 0.00740196
R1569 iovss.n680 iovss.n679 0.00740196
R1570 iovss.n739 iovss 0.00727871
R1571 iovss.n1016 iovss.n2 0.00727735
R1572 iovss.n1019 iovss.n1018 0.00716247
R1573 iovss.n160 iovss 0.00671176
R1574 iovss.n774 iovss.n1 0.00666247
R1575 iovss.n778 iovss.n1 0.00627731
R1576 iovss.n5 iovss.n1 0.0057381
R1577 iovss.n775 iovss.n1 0.0057381
R1578 iovss.n444 iovss.n1 0.00565631
R1579 iovss.n873 iovss.n872 0.0047102
R1580 iovss.n899 iovss.n113 0.0047102
R1581 iovss.n240 iovss.n239 0.00442211
R1582 iovss.n547 iovss.n546 0.00442211
R1583 iovss.n242 iovss.n241 0.00395098
R1584 iovss.n245 iovss.n241 0.00395098
R1585 iovss.n247 iovss.n245 0.00395098
R1586 iovss.n247 iovss.n246 0.00395098
R1587 iovss.n246 iovss.n236 0.00395098
R1588 iovss.n254 iovss.n236 0.00395098
R1589 iovss.n254 iovss.n253 0.00395098
R1590 iovss.n253 iovss.n237 0.00395098
R1591 iovss.n237 iovss.n232 0.00395098
R1592 iovss.n260 iovss.n232 0.00395098
R1593 iovss.n262 iovss.n260 0.00395098
R1594 iovss.n262 iovss.n261 0.00395098
R1595 iovss.n261 iovss.n227 0.00395098
R1596 iovss.n269 iovss.n227 0.00395098
R1597 iovss.n269 iovss.n268 0.00395098
R1598 iovss.n268 iovss.n228 0.00395098
R1599 iovss.n228 iovss.n223 0.00395098
R1600 iovss.n275 iovss.n223 0.00395098
R1601 iovss.n277 iovss.n275 0.00395098
R1602 iovss.n277 iovss.n276 0.00395098
R1603 iovss.n276 iovss.n218 0.00395098
R1604 iovss.n284 iovss.n218 0.00395098
R1605 iovss.n284 iovss.n283 0.00395098
R1606 iovss.n283 iovss.n219 0.00395098
R1607 iovss.n219 iovss.n214 0.00395098
R1608 iovss.n290 iovss.n214 0.00395098
R1609 iovss.n292 iovss.n290 0.00395098
R1610 iovss.n292 iovss.n291 0.00395098
R1611 iovss.n291 iovss.n209 0.00395098
R1612 iovss.n299 iovss.n209 0.00395098
R1613 iovss.n299 iovss.n298 0.00395098
R1614 iovss.n298 iovss.n210 0.00395098
R1615 iovss.n210 iovss.n205 0.00395098
R1616 iovss.n305 iovss.n205 0.00395098
R1617 iovss.n307 iovss.n305 0.00395098
R1618 iovss.n307 iovss.n306 0.00395098
R1619 iovss.n306 iovss.n200 0.00395098
R1620 iovss.n314 iovss.n200 0.00395098
R1621 iovss.n314 iovss.n313 0.00395098
R1622 iovss.n313 iovss.n201 0.00395098
R1623 iovss.n201 iovss.n196 0.00395098
R1624 iovss.n320 iovss.n196 0.00395098
R1625 iovss.n322 iovss.n320 0.00395098
R1626 iovss.n322 iovss.n321 0.00395098
R1627 iovss.n321 iovss.n191 0.00395098
R1628 iovss.n329 iovss.n191 0.00395098
R1629 iovss.n329 iovss.n328 0.00395098
R1630 iovss.n328 iovss.n192 0.00395098
R1631 iovss.n192 iovss.n187 0.00395098
R1632 iovss.n335 iovss.n187 0.00395098
R1633 iovss.n337 iovss.n335 0.00395098
R1634 iovss.n337 iovss.n336 0.00395098
R1635 iovss.n336 iovss.n182 0.00395098
R1636 iovss.n344 iovss.n182 0.00395098
R1637 iovss.n344 iovss.n343 0.00395098
R1638 iovss.n343 iovss.n183 0.00395098
R1639 iovss.n183 iovss.n178 0.00395098
R1640 iovss.n350 iovss.n178 0.00395098
R1641 iovss.n352 iovss.n350 0.00395098
R1642 iovss.n352 iovss.n351 0.00395098
R1643 iovss.n351 iovss.n173 0.00395098
R1644 iovss.n359 iovss.n173 0.00395098
R1645 iovss.n359 iovss.n358 0.00395098
R1646 iovss.n358 iovss.n174 0.00395098
R1647 iovss.n174 iovss.n169 0.00395098
R1648 iovss.n365 iovss.n169 0.00395098
R1649 iovss.n367 iovss.n365 0.00395098
R1650 iovss.n367 iovss.n366 0.00395098
R1651 iovss.n366 iovss.n166 0.00395098
R1652 iovss.n877 iovss.n166 0.00395098
R1653 iovss.n877 iovss.n876 0.00395098
R1654 iovss.n876 iovss.n167 0.00395098
R1655 iovss.n167 iovss.n162 0.00395098
R1656 iovss.n883 iovss.n162 0.00395098
R1657 iovss.n548 iovss.n545 0.00395098
R1658 iovss.n550 iovss.n548 0.00395098
R1659 iovss.n550 iovss.n549 0.00395098
R1660 iovss.n549 iovss.n542 0.00395098
R1661 iovss.n557 iovss.n542 0.00395098
R1662 iovss.n557 iovss.n556 0.00395098
R1663 iovss.n556 iovss.n543 0.00395098
R1664 iovss.n543 iovss.n538 0.00395098
R1665 iovss.n563 iovss.n538 0.00395098
R1666 iovss.n565 iovss.n563 0.00395098
R1667 iovss.n565 iovss.n564 0.00395098
R1668 iovss.n564 iovss.n533 0.00395098
R1669 iovss.n572 iovss.n533 0.00395098
R1670 iovss.n572 iovss.n571 0.00395098
R1671 iovss.n571 iovss.n534 0.00395098
R1672 iovss.n534 iovss.n529 0.00395098
R1673 iovss.n578 iovss.n529 0.00395098
R1674 iovss.n580 iovss.n578 0.00395098
R1675 iovss.n580 iovss.n579 0.00395098
R1676 iovss.n579 iovss.n524 0.00395098
R1677 iovss.n587 iovss.n524 0.00395098
R1678 iovss.n587 iovss.n586 0.00395098
R1679 iovss.n586 iovss.n525 0.00395098
R1680 iovss.n525 iovss.n520 0.00395098
R1681 iovss.n593 iovss.n520 0.00395098
R1682 iovss.n595 iovss.n593 0.00395098
R1683 iovss.n595 iovss.n594 0.00395098
R1684 iovss.n594 iovss.n515 0.00395098
R1685 iovss.n602 iovss.n515 0.00395098
R1686 iovss.n602 iovss.n601 0.00395098
R1687 iovss.n601 iovss.n516 0.00395098
R1688 iovss.n516 iovss.n511 0.00395098
R1689 iovss.n608 iovss.n511 0.00395098
R1690 iovss.n610 iovss.n608 0.00395098
R1691 iovss.n610 iovss.n609 0.00395098
R1692 iovss.n609 iovss.n506 0.00395098
R1693 iovss.n617 iovss.n506 0.00395098
R1694 iovss.n617 iovss.n616 0.00395098
R1695 iovss.n616 iovss.n507 0.00395098
R1696 iovss.n507 iovss.n502 0.00395098
R1697 iovss.n623 iovss.n502 0.00395098
R1698 iovss.n625 iovss.n623 0.00395098
R1699 iovss.n625 iovss.n624 0.00395098
R1700 iovss.n624 iovss.n497 0.00395098
R1701 iovss.n632 iovss.n497 0.00395098
R1702 iovss.n632 iovss.n631 0.00395098
R1703 iovss.n631 iovss.n498 0.00395098
R1704 iovss.n498 iovss.n493 0.00395098
R1705 iovss.n638 iovss.n493 0.00395098
R1706 iovss.n640 iovss.n638 0.00395098
R1707 iovss.n640 iovss.n639 0.00395098
R1708 iovss.n639 iovss.n488 0.00395098
R1709 iovss.n647 iovss.n488 0.00395098
R1710 iovss.n647 iovss.n646 0.00395098
R1711 iovss.n646 iovss.n489 0.00395098
R1712 iovss.n489 iovss.n484 0.00395098
R1713 iovss.n653 iovss.n484 0.00395098
R1714 iovss.n655 iovss.n653 0.00395098
R1715 iovss.n655 iovss.n654 0.00395098
R1716 iovss.n654 iovss.n479 0.00395098
R1717 iovss.n662 iovss.n479 0.00395098
R1718 iovss.n662 iovss.n661 0.00395098
R1719 iovss.n661 iovss.n480 0.00395098
R1720 iovss.n480 iovss.n475 0.00395098
R1721 iovss.n668 iovss.n475 0.00395098
R1722 iovss.n670 iovss.n668 0.00395098
R1723 iovss.n670 iovss.n669 0.00395098
R1724 iovss.n669 iovss.n470 0.00395098
R1725 iovss.n686 iovss.n470 0.00395098
R1726 iovss.n686 iovss.n685 0.00395098
R1727 iovss.n685 iovss.n471 0.00395098
R1728 iovss.n682 iovss.n471 0.00395098
R1729 iovss.n682 iovss.n681 0.00395098
R1730 iovss.n681 iovss.n678 0.00395098
R1731 iovss iovss.n1020 0.00358123
R1732 iovss.n1001 iovss.n57 0.00326078
R1733 iovss.n906 iovss.n72 0.00326078
R1734 iovss.n745 iovss.n740 0.00314333
R1735 iovss.n697 iovss.n1 0.00306909
R1736 iovss.n742 iovss.n741 0.00298471
R1737 iovss.n692 iovss.n688 0.00298471
R1738 iovss.n445 iovss.n444 0.00261959
R1739 iovss.n677 iovss 0.00261765
R1740 iovss.n442 iovss.n0 0.00248367
R1741 iovss.n66 iovss.n65 0.00219098
R1742 iovss.n906 iovss.n66 0.00219098
R1743 iovss.n1019 iovss.n2 0.00199991
R1744 iovss.n676 iovss 0.00196667
R1745 iovss.n881 iovss 0.00196667
R1746 iovss.n244 iovss.n235 0.00191176
R1747 iovss.n255 iovss.n235 0.00191176
R1748 iovss.n255 iovss.n233 0.00191176
R1749 iovss.n259 iovss.n233 0.00191176
R1750 iovss.n259 iovss.n226 0.00191176
R1751 iovss.n270 iovss.n226 0.00191176
R1752 iovss.n270 iovss.n224 0.00191176
R1753 iovss.n274 iovss.n224 0.00191176
R1754 iovss.n274 iovss.n217 0.00191176
R1755 iovss.n285 iovss.n217 0.00191176
R1756 iovss.n285 iovss.n215 0.00191176
R1757 iovss.n289 iovss.n215 0.00191176
R1758 iovss.n289 iovss.n208 0.00191176
R1759 iovss.n300 iovss.n208 0.00191176
R1760 iovss.n300 iovss.n206 0.00191176
R1761 iovss.n304 iovss.n206 0.00191176
R1762 iovss.n304 iovss.n199 0.00191176
R1763 iovss.n315 iovss.n199 0.00191176
R1764 iovss.n315 iovss.n197 0.00191176
R1765 iovss.n319 iovss.n197 0.00191176
R1766 iovss.n319 iovss.n190 0.00191176
R1767 iovss.n330 iovss.n190 0.00191176
R1768 iovss.n330 iovss.n188 0.00191176
R1769 iovss.n334 iovss.n188 0.00191176
R1770 iovss.n334 iovss.n181 0.00191176
R1771 iovss.n345 iovss.n181 0.00191176
R1772 iovss.n345 iovss.n179 0.00191176
R1773 iovss.n349 iovss.n179 0.00191176
R1774 iovss.n349 iovss.n172 0.00191176
R1775 iovss.n360 iovss.n172 0.00191176
R1776 iovss.n360 iovss.n170 0.00191176
R1777 iovss.n364 iovss.n170 0.00191176
R1778 iovss.n364 iovss.n165 0.00191176
R1779 iovss.n878 iovss.n165 0.00191176
R1780 iovss.n878 iovss.n163 0.00191176
R1781 iovss.n882 iovss.n163 0.00191176
R1782 iovss.n551 iovss.n544 0.00191176
R1783 iovss.n555 iovss.n544 0.00191176
R1784 iovss.n555 iovss.n537 0.00191176
R1785 iovss.n566 iovss.n537 0.00191176
R1786 iovss.n566 iovss.n535 0.00191176
R1787 iovss.n570 iovss.n535 0.00191176
R1788 iovss.n570 iovss.n528 0.00191176
R1789 iovss.n581 iovss.n528 0.00191176
R1790 iovss.n581 iovss.n526 0.00191176
R1791 iovss.n585 iovss.n526 0.00191176
R1792 iovss.n585 iovss.n519 0.00191176
R1793 iovss.n596 iovss.n519 0.00191176
R1794 iovss.n596 iovss.n517 0.00191176
R1795 iovss.n600 iovss.n517 0.00191176
R1796 iovss.n600 iovss.n510 0.00191176
R1797 iovss.n611 iovss.n510 0.00191176
R1798 iovss.n611 iovss.n508 0.00191176
R1799 iovss.n615 iovss.n508 0.00191176
R1800 iovss.n615 iovss.n501 0.00191176
R1801 iovss.n626 iovss.n501 0.00191176
R1802 iovss.n626 iovss.n499 0.00191176
R1803 iovss.n630 iovss.n499 0.00191176
R1804 iovss.n630 iovss.n492 0.00191176
R1805 iovss.n641 iovss.n492 0.00191176
R1806 iovss.n641 iovss.n490 0.00191176
R1807 iovss.n645 iovss.n490 0.00191176
R1808 iovss.n645 iovss.n483 0.00191176
R1809 iovss.n656 iovss.n483 0.00191176
R1810 iovss.n656 iovss.n481 0.00191176
R1811 iovss.n660 iovss.n481 0.00191176
R1812 iovss.n660 iovss.n474 0.00191176
R1813 iovss.n671 iovss.n474 0.00191176
R1814 iovss.n671 iovss.n472 0.00191176
R1815 iovss.n684 iovss.n472 0.00191176
R1816 iovss.n684 iovss.n683 0.00191176
R1817 iovss.n683 iovss.n677 0.00191176
R1818 iovss.n893 iovss.n96 0.00189683
R1819 iovss.n887 iovss.n886 0.00189683
R1820 iovss.n703 iovss.n448 0.00189683
R1821 iovss.n736 iovss.n711 0.00189683
R1822 iovss.n66 iovss.n61 0.00189683
R1823 iovss.n914 iovss.n10 0.00189683
R1824 iovss.n1012 iovss.n10 0.00184541
R1825 iovss.n1001 iovss.n6 0.00184541
R1826 iovss.n737 iovss.n736 0.00184541
R1827 iovss.n747 iovss.n370 0.00184541
R1828 iovss.n886 iovss.n134 0.00184541
R1829 iovss.n1012 iovss.n1011 0.00184541
R1830 iovss.n10 iovss.n6 0.00184541
R1831 iovss.n736 iovss.n370 0.00184541
R1832 iovss.n742 iovss.n737 0.00184541
R1833 iovss.n872 iovss.n134 0.00184541
R1834 iovss.n450 iovss.n448 0.00184541
R1835 iovss.n464 iovss.n448 0.00184541
R1836 iovss.n117 iovss.n96 0.00184541
R1837 iovss.n899 iovss.n117 0.00184541
R1838 iovss.n692 iovss.n450 0.00184541
R1839 iovss.n699 iovss.n464 0.00184541
R1840 iovss.n697 iovss.n696 0.00171968
R1841 iovss.n244 iovss.n243 0.0016983
R1842 iovss.n552 iovss.n551 0.0016983
R1843 iovss.n874 iovss.n747 0.00153529
R1844 iovss.n699 iovss.n458 0.00153529
R1845 iovss.n886 iovss.n885 0.00150078
R1846 iovss.n98 iovss.n96 0.00150078
R1847 iovss.n740 iovss.n1 0.00149998
R1848 iovss.n740 iovss.n739 0.00149998
R1849 iovss.n442 iovss.n1 0.00149997
R1850 iovss.n2 iovss.n1 0.00149991
R1851 iovss.n738 iovss.n1 0.0014837
R1852 iovss.n1020 iovss.n0 0.0014837
R1853 iovss.n739 iovss.n738 0.0014837
R1854 iovss.n554 iovss.n553 0.00147778
R1855 iovss.n554 iovss.n536 0.00147778
R1856 iovss.n567 iovss.n536 0.00147778
R1857 iovss.n568 iovss.n567 0.00147778
R1858 iovss.n569 iovss.n568 0.00147778
R1859 iovss.n569 iovss.n527 0.00147778
R1860 iovss.n582 iovss.n527 0.00147778
R1861 iovss.n583 iovss.n582 0.00147778
R1862 iovss.n584 iovss.n583 0.00147778
R1863 iovss.n584 iovss.n518 0.00147778
R1864 iovss.n597 iovss.n518 0.00147778
R1865 iovss.n598 iovss.n597 0.00147778
R1866 iovss.n599 iovss.n598 0.00147778
R1867 iovss.n599 iovss.n509 0.00147778
R1868 iovss.n612 iovss.n509 0.00147778
R1869 iovss.n613 iovss.n612 0.00147778
R1870 iovss.n614 iovss.n613 0.00147778
R1871 iovss.n614 iovss.n500 0.00147778
R1872 iovss.n627 iovss.n500 0.00147778
R1873 iovss.n628 iovss.n627 0.00147778
R1874 iovss.n629 iovss.n628 0.00147778
R1875 iovss.n629 iovss.n491 0.00147778
R1876 iovss.n642 iovss.n491 0.00147778
R1877 iovss.n643 iovss.n642 0.00147778
R1878 iovss.n644 iovss.n643 0.00147778
R1879 iovss.n644 iovss.n482 0.00147778
R1880 iovss.n657 iovss.n482 0.00147778
R1881 iovss.n658 iovss.n657 0.00147778
R1882 iovss.n659 iovss.n658 0.00147778
R1883 iovss.n659 iovss.n473 0.00147778
R1884 iovss.n672 iovss.n473 0.00147778
R1885 iovss.n673 iovss.n672 0.00147778
R1886 iovss.n674 iovss.n673 0.00147778
R1887 iovss.n675 iovss.n674 0.00147778
R1888 iovss.n676 iovss.n675 0.00147778
R1889 iovss.n256 iovss.n234 0.00147778
R1890 iovss.n257 iovss.n256 0.00147778
R1891 iovss.n258 iovss.n257 0.00147778
R1892 iovss.n258 iovss.n225 0.00147778
R1893 iovss.n271 iovss.n225 0.00147778
R1894 iovss.n272 iovss.n271 0.00147778
R1895 iovss.n273 iovss.n272 0.00147778
R1896 iovss.n273 iovss.n216 0.00147778
R1897 iovss.n286 iovss.n216 0.00147778
R1898 iovss.n287 iovss.n286 0.00147778
R1899 iovss.n288 iovss.n287 0.00147778
R1900 iovss.n288 iovss.n207 0.00147778
R1901 iovss.n301 iovss.n207 0.00147778
R1902 iovss.n302 iovss.n301 0.00147778
R1903 iovss.n303 iovss.n302 0.00147778
R1904 iovss.n303 iovss.n198 0.00147778
R1905 iovss.n316 iovss.n198 0.00147778
R1906 iovss.n317 iovss.n316 0.00147778
R1907 iovss.n318 iovss.n317 0.00147778
R1908 iovss.n318 iovss.n189 0.00147778
R1909 iovss.n331 iovss.n189 0.00147778
R1910 iovss.n332 iovss.n331 0.00147778
R1911 iovss.n333 iovss.n332 0.00147778
R1912 iovss.n333 iovss.n180 0.00147778
R1913 iovss.n346 iovss.n180 0.00147778
R1914 iovss.n347 iovss.n346 0.00147778
R1915 iovss.n348 iovss.n347 0.00147778
R1916 iovss.n348 iovss.n171 0.00147778
R1917 iovss.n361 iovss.n171 0.00147778
R1918 iovss.n362 iovss.n361 0.00147778
R1919 iovss.n363 iovss.n362 0.00147778
R1920 iovss.n363 iovss.n164 0.00147778
R1921 iovss.n879 iovss.n164 0.00147778
R1922 iovss.n880 iovss.n879 0.00147778
R1923 iovss.n881 iovss.n880 0.00147778
R1924 iovss.n452 iovss.n1 0.00133247
R1925 iovss.n1011 iovss.n11 0.00125922
R1926 iovss.n666 iovss.n65 0.00125922
R1927 iovss.n885 iovss.n160 0.0011902
R1928 iovss.n902 iovss.n98 0.0011902
R1929 iovss.n904 iovss.n1 0.00109598
R1930 iovss.n1020 iovss.n1019 0.001
R1931 iovdd.n1307 iovdd.n43 17.0005
R1932 iovdd.n1307 iovdd.n5 17.0005
R1933 iovdd.n49 iovdd.n43 17.0005
R1934 iovdd.n49 iovdd.n4 17.0005
R1935 iovdd.n1359 iovdd.n49 17.0005
R1936 iovdd.n49 iovdd.n42 17.0005
R1937 iovdd.n49 iovdd.n40 17.0005
R1938 iovdd.n49 iovdd.n39 17.0005
R1939 iovdd.n49 iovdd.n37 17.0005
R1940 iovdd.n49 iovdd.n36 17.0005
R1941 iovdd.n49 iovdd.n34 17.0005
R1942 iovdd.n49 iovdd.n33 17.0005
R1943 iovdd.n49 iovdd.n31 17.0005
R1944 iovdd.n49 iovdd.n30 17.0005
R1945 iovdd.n49 iovdd.n28 17.0005
R1946 iovdd.n49 iovdd.n27 17.0005
R1947 iovdd.n49 iovdd.n23 17.0005
R1948 iovdd.n49 iovdd.n22 17.0005
R1949 iovdd.n49 iovdd.n20 17.0005
R1950 iovdd.n49 iovdd.n19 17.0005
R1951 iovdd.n49 iovdd.n17 17.0005
R1952 iovdd.n49 iovdd.n16 17.0005
R1953 iovdd.n49 iovdd.n13 17.0005
R1954 iovdd.n49 iovdd.n12 17.0005
R1955 iovdd.n49 iovdd.n11 17.0005
R1956 iovdd.n49 iovdd.n10 17.0005
R1957 iovdd.n49 iovdd.n9 17.0005
R1958 iovdd.n1229 iovdd.n49 17.0005
R1959 iovdd.n49 iovdd.n7 17.0005
R1960 iovdd.n49 iovdd.n5 17.0005
R1961 iovdd.n1313 iovdd.n272 9.0005
R1962 iovdd.n1313 iovdd.n273 9.0005
R1963 iovdd.n547 iovdd.n479 9.0005
R1964 iovdd.n547 iovdd.n483 9.0005
R1965 iovdd.n547 iovdd.n476 9.0005
R1966 iovdd.n547 iovdd.n486 9.0005
R1967 iovdd.n547 iovdd.n474 9.0005
R1968 iovdd.n547 iovdd.n489 9.0005
R1969 iovdd.n547 iovdd.n472 9.0005
R1970 iovdd.n547 iovdd.n492 9.0005
R1971 iovdd.n547 iovdd.n470 9.0005
R1972 iovdd.n547 iovdd.n495 9.0005
R1973 iovdd.n547 iovdd.n468 9.0005
R1974 iovdd.n547 iovdd.n498 9.0005
R1975 iovdd.n547 iovdd.n466 9.0005
R1976 iovdd.n547 iovdd.n501 9.0005
R1977 iovdd.n547 iovdd.n464 9.0005
R1978 iovdd.n547 iovdd.n504 9.0005
R1979 iovdd.n547 iovdd.n462 9.0005
R1980 iovdd.n547 iovdd.n507 9.0005
R1981 iovdd.n547 iovdd.n460 9.0005
R1982 iovdd.n547 iovdd.n510 9.0005
R1983 iovdd.n547 iovdd.n458 9.0005
R1984 iovdd.n547 iovdd.n513 9.0005
R1985 iovdd.n547 iovdd.n456 9.0005
R1986 iovdd.n547 iovdd.n516 9.0005
R1987 iovdd.n547 iovdd.n454 9.0005
R1988 iovdd.n547 iovdd.n519 9.0005
R1989 iovdd.n547 iovdd.n452 9.0005
R1990 iovdd.n547 iovdd.n522 9.0005
R1991 iovdd.n547 iovdd.n450 9.0005
R1992 iovdd.n547 iovdd.n525 9.0005
R1993 iovdd.n547 iovdd.n448 9.0005
R1994 iovdd.n547 iovdd.n528 9.0005
R1995 iovdd.n547 iovdd.n446 9.0005
R1996 iovdd.n547 iovdd.n531 9.0005
R1997 iovdd.n547 iovdd.n444 9.0005
R1998 iovdd.n547 iovdd.n534 9.0005
R1999 iovdd.n547 iovdd.n442 9.0005
R2000 iovdd.n547 iovdd.n537 9.0005
R2001 iovdd.n547 iovdd.n440 9.0005
R2002 iovdd.n547 iovdd.n540 9.0005
R2003 iovdd.n547 iovdd.n438 9.0005
R2004 iovdd.n547 iovdd.n543 9.0005
R2005 iovdd.n547 iovdd.n436 9.0005
R2006 iovdd.n547 iovdd.n546 9.0005
R2007 iovdd.n547 iovdd.n434 9.0005
R2008 iovdd.n1313 iovdd.n1312 9.0005
R2009 iovdd.n1223 iovdd.n862 9.0005
R2010 iovdd.n1221 iovdd.n862 9.0005
R2011 iovdd.n1218 iovdd.n862 9.0005
R2012 iovdd.n1221 iovdd.n1136 9.0005
R2013 iovdd.n1221 iovdd.n1138 9.0005
R2014 iovdd.n1221 iovdd.n1134 9.0005
R2015 iovdd.n1221 iovdd.n1140 9.0005
R2016 iovdd.n1221 iovdd.n1132 9.0005
R2017 iovdd.n1221 iovdd.n1142 9.0005
R2018 iovdd.n1221 iovdd.n1130 9.0005
R2019 iovdd.n1221 iovdd.n1144 9.0005
R2020 iovdd.n1221 iovdd.n1128 9.0005
R2021 iovdd.n1221 iovdd.n1146 9.0005
R2022 iovdd.n1221 iovdd.n1126 9.0005
R2023 iovdd.n1221 iovdd.n1148 9.0005
R2024 iovdd.n1221 iovdd.n1124 9.0005
R2025 iovdd.n1221 iovdd.n1150 9.0005
R2026 iovdd.n1221 iovdd.n1122 9.0005
R2027 iovdd.n1221 iovdd.n1152 9.0005
R2028 iovdd.n1221 iovdd.n1120 9.0005
R2029 iovdd.n1221 iovdd.n1154 9.0005
R2030 iovdd.n1221 iovdd.n1118 9.0005
R2031 iovdd.n1221 iovdd.n1156 9.0005
R2032 iovdd.n1221 iovdd.n1116 9.0005
R2033 iovdd.n1221 iovdd.n1158 9.0005
R2034 iovdd.n1221 iovdd.n1114 9.0005
R2035 iovdd.n1221 iovdd.n1160 9.0005
R2036 iovdd.n1221 iovdd.n1112 9.0005
R2037 iovdd.n1221 iovdd.n1162 9.0005
R2038 iovdd.n1221 iovdd.n1110 9.0005
R2039 iovdd.n1221 iovdd.n1164 9.0005
R2040 iovdd.n1221 iovdd.n1108 9.0005
R2041 iovdd.n1221 iovdd.n1166 9.0005
R2042 iovdd.n1221 iovdd.n1106 9.0005
R2043 iovdd.n1221 iovdd.n1168 9.0005
R2044 iovdd.n1221 iovdd.n1104 9.0005
R2045 iovdd.n1221 iovdd.n1170 9.0005
R2046 iovdd.n1221 iovdd.n1102 9.0005
R2047 iovdd.n1221 iovdd.n1172 9.0005
R2048 iovdd.n1221 iovdd.n1100 9.0005
R2049 iovdd.n1221 iovdd.n1174 9.0005
R2050 iovdd.n1221 iovdd.n1098 9.0005
R2051 iovdd.n1221 iovdd.n1176 9.0005
R2052 iovdd.n1221 iovdd.n1096 9.0005
R2053 iovdd.n1221 iovdd.n1178 9.0005
R2054 iovdd.n1221 iovdd.n1094 9.0005
R2055 iovdd.n1221 iovdd.n1180 9.0005
R2056 iovdd.n1221 iovdd.n1092 9.0005
R2057 iovdd.n1221 iovdd.n1220 9.0005
R2058 iovdd.n1220 iovdd.n1218 9.0005
R2059 iovdd.n1218 iovdd.n860 9.0005
R2060 iovdd.n1221 iovdd.n860 9.0005
R2061 iovdd.n297 iovdd.n290 9.0005
R2062 iovdd.n297 iovdd.n275 9.0005
R2063 iovdd.n1311 iovdd.n297 9.0005
R2064 iovdd.n1225 iovdd.n860 9.0005
R2065 iovdd.n1227 iovdd.n860 9.0005
R2066 iovdd.n863 iovdd.n860 9.0005
R2067 iovdd.n1312 iovdd.n290 9.0005
R2068 iovdd.n1312 iovdd.n275 9.0005
R2069 iovdd.n1312 iovdd.n1311 9.0005
R2070 iovdd.n1226 iovdd.n1225 9.0005
R2071 iovdd.n1226 iovdd.n863 9.0005
R2072 iovdd.n1227 iovdd.n1226 9.0005
R2073 iovdd.n1357 iovdd.n113 9.0005
R2074 iovdd.n113 iovdd.n111 9.0005
R2075 iovdd.n1357 iovdd.n1356 9.0005
R2076 iovdd.n1355 iovdd.n165 9.0005
R2077 iovdd.n1355 iovdd.n168 9.0005
R2078 iovdd.n1355 iovdd.n164 9.0005
R2079 iovdd.n1355 iovdd.n171 9.0005
R2080 iovdd.n1355 iovdd.n162 9.0005
R2081 iovdd.n1355 iovdd.n174 9.0005
R2082 iovdd.n1355 iovdd.n160 9.0005
R2083 iovdd.n1355 iovdd.n177 9.0005
R2084 iovdd.n1355 iovdd.n158 9.0005
R2085 iovdd.n1355 iovdd.n180 9.0005
R2086 iovdd.n1355 iovdd.n156 9.0005
R2087 iovdd.n1355 iovdd.n183 9.0005
R2088 iovdd.n1355 iovdd.n154 9.0005
R2089 iovdd.n1355 iovdd.n186 9.0005
R2090 iovdd.n1355 iovdd.n152 9.0005
R2091 iovdd.n1355 iovdd.n189 9.0005
R2092 iovdd.n1355 iovdd.n150 9.0005
R2093 iovdd.n1355 iovdd.n192 9.0005
R2094 iovdd.n1355 iovdd.n148 9.0005
R2095 iovdd.n1355 iovdd.n195 9.0005
R2096 iovdd.n1355 iovdd.n146 9.0005
R2097 iovdd.n1355 iovdd.n198 9.0005
R2098 iovdd.n1355 iovdd.n144 9.0005
R2099 iovdd.n1355 iovdd.n201 9.0005
R2100 iovdd.n1355 iovdd.n142 9.0005
R2101 iovdd.n1355 iovdd.n204 9.0005
R2102 iovdd.n1355 iovdd.n140 9.0005
R2103 iovdd.n1355 iovdd.n207 9.0005
R2104 iovdd.n1355 iovdd.n138 9.0005
R2105 iovdd.n1355 iovdd.n210 9.0005
R2106 iovdd.n1355 iovdd.n136 9.0005
R2107 iovdd.n1355 iovdd.n213 9.0005
R2108 iovdd.n1355 iovdd.n134 9.0005
R2109 iovdd.n1355 iovdd.n216 9.0005
R2110 iovdd.n1355 iovdd.n132 9.0005
R2111 iovdd.n1355 iovdd.n219 9.0005
R2112 iovdd.n1355 iovdd.n130 9.0005
R2113 iovdd.n1355 iovdd.n222 9.0005
R2114 iovdd.n1355 iovdd.n128 9.0005
R2115 iovdd.n1355 iovdd.n225 9.0005
R2116 iovdd.n1355 iovdd.n126 9.0005
R2117 iovdd.n1355 iovdd.n228 9.0005
R2118 iovdd.n1355 iovdd.n124 9.0005
R2119 iovdd.n1355 iovdd.n231 9.0005
R2120 iovdd.n1355 iovdd.n122 9.0005
R2121 iovdd.n1355 iovdd.n234 9.0005
R2122 iovdd.n1355 iovdd.n120 9.0005
R2123 iovdd.n1354 iovdd.n1353 9.0005
R2124 iovdd.n1355 iovdd.n1354 9.0005
R2125 iovdd.n1356 iovdd.n115 9.0005
R2126 iovdd.n1356 iovdd.n1355 9.0005
R2127 iovdd.n1355 iovdd.n113 9.0005
R2128 iovdd.n1356 iovdd.n111 9.0005
R2129 iovdd.n1301 iovdd.n1300 9.0005
R2130 iovdd.n1304 iovdd.n400 9.0005
R2131 iovdd.n1304 iovdd.n404 9.0005
R2132 iovdd.n1304 iovdd.n398 9.0005
R2133 iovdd.n1304 iovdd.n407 9.0005
R2134 iovdd.n1304 iovdd.n396 9.0005
R2135 iovdd.n1304 iovdd.n410 9.0005
R2136 iovdd.n1304 iovdd.n394 9.0005
R2137 iovdd.n1304 iovdd.n1303 9.0005
R2138 iovdd.n1304 iovdd.n392 9.0005
R2139 iovdd.n1305 iovdd.n389 9.0005
R2140 iovdd.n1305 iovdd.n1304 9.0005
R2141 iovdd.n1264 iovdd.n424 9.0005
R2142 iovdd.n1261 iovdd.n424 9.0005
R2143 iovdd.n1261 iovdd.n1251 9.0005
R2144 iovdd.n1261 iovdd.n1248 9.0005
R2145 iovdd.n1261 iovdd.n1254 9.0005
R2146 iovdd.n1261 iovdd.n1246 9.0005
R2147 iovdd.n1261 iovdd.n1257 9.0005
R2148 iovdd.n1261 iovdd.n1244 9.0005
R2149 iovdd.n1261 iovdd.n1260 9.0005
R2150 iovdd.n1261 iovdd.n1242 9.0005
R2151 iovdd.n1262 iovdd.n1261 9.0005
R2152 iovdd.n1261 iovdd.n565 9.0005
R2153 iovdd.n1264 iovdd.n388 9.0005
R2154 iovdd.n1261 iovdd.n388 9.0005
R2155 iovdd.n1236 iovdd.n771 9.0005
R2156 iovdd.n1233 iovdd.n771 9.0005
R2157 iovdd.n1233 iovdd.n786 9.0005
R2158 iovdd.n1233 iovdd.n784 9.0005
R2159 iovdd.n1233 iovdd.n788 9.0005
R2160 iovdd.n1233 iovdd.n783 9.0005
R2161 iovdd.n1233 iovdd.n1232 9.0005
R2162 iovdd.n1233 iovdd.n782 9.0005
R2163 iovdd.n1234 iovdd.n1233 9.0005
R2164 iovdd.n1233 iovdd.n778 9.0005
R2165 iovdd.n1237 iovdd.n1236 9.0005
R2166 iovdd.n774 iovdd.n773 9.0005
R2167 iovdd.n1307 iovdd.n47 8.501
R2168 iovdd.n1307 iovdd.n386 8.501
R2169 iovdd.n1307 iovdd.n385 8.501
R2170 iovdd.n1307 iovdd.n384 8.501
R2171 iovdd.n1307 iovdd.n383 8.501
R2172 iovdd.n1307 iovdd.n382 8.501
R2173 iovdd.n1307 iovdd.n362 8.501
R2174 iovdd.n1308 iovdd.n1307 8.501
R2175 iovdd.n1307 iovdd.n381 8.501
R2176 iovdd.n1307 iovdd.n380 8.501
R2177 iovdd.n1307 iovdd.n379 8.501
R2178 iovdd.n1307 iovdd.n378 8.501
R2179 iovdd.n1307 iovdd.n377 8.501
R2180 iovdd.n1307 iovdd.n376 8.501
R2181 iovdd.n375 iovdd.n374 8.501
R2182 iovdd.n375 iovdd.n48 8.501
R2183 iovdd.n375 iovdd.n373 8.501
R2184 iovdd.n375 iovdd.n372 8.501
R2185 iovdd.n375 iovdd.n371 8.501
R2186 iovdd.n375 iovdd.n370 8.501
R2187 iovdd.n375 iovdd.n369 8.501
R2188 iovdd.n375 iovdd.n368 8.501
R2189 iovdd.n375 iovdd.n367 8.501
R2190 iovdd.n375 iovdd.n366 8.501
R2191 iovdd.n375 iovdd.n365 8.501
R2192 iovdd.n375 iovdd.n364 8.501
R2193 iovdd.n857 iovdd.n375 8.501
R2194 iovdd.n375 iovdd.n363 8.501
R2195 iovdd.n1309 iovdd.n375 8.5005
R2196 iovdd.n1309 iovdd.n49 8.5005
R2197 iovdd.n1360 iovdd.n44 5.66866
R2198 iovdd.n858 iovdd.n6 5.66767
R2199 iovdd.n1309 iovdd.n359 5.66717
R2200 iovdd.n1309 iovdd.n357 5.66717
R2201 iovdd.n1309 iovdd.n356 5.66717
R2202 iovdd.n1309 iovdd.n354 5.66717
R2203 iovdd.n1309 iovdd.n352 5.66717
R2204 iovdd.n1309 iovdd.n350 5.66717
R2205 iovdd.n1309 iovdd.n348 5.66717
R2206 iovdd.n1309 iovdd.n347 5.66717
R2207 iovdd.n1309 iovdd.n345 5.66717
R2208 iovdd.n1309 iovdd.n343 5.66717
R2209 iovdd.n1309 iovdd.n341 5.66717
R2210 iovdd.n1309 iovdd.n339 5.66717
R2211 iovdd.n1309 iovdd.n338 5.66717
R2212 iovdd.n1309 iovdd.n336 5.66717
R2213 iovdd.n1309 iovdd.n334 5.66717
R2214 iovdd.n1309 iovdd.n332 5.66717
R2215 iovdd.n1309 iovdd.n330 5.66717
R2216 iovdd.n1309 iovdd.n329 5.66717
R2217 iovdd.n1309 iovdd.n327 5.66717
R2218 iovdd.n1309 iovdd.n325 5.66717
R2219 iovdd.n1309 iovdd.n323 5.66717
R2220 iovdd.n1309 iovdd.n322 5.66717
R2221 iovdd.n1309 iovdd.n320 5.66717
R2222 iovdd.n1309 iovdd.n318 5.66717
R2223 iovdd.n1309 iovdd.n316 5.66717
R2224 iovdd.n1309 iovdd.n314 5.66717
R2225 iovdd.n1309 iovdd.n313 5.66717
R2226 iovdd.n1309 iovdd.n311 5.66717
R2227 iovdd.n1309 iovdd.n309 5.66717
R2228 iovdd.n1309 iovdd.n307 5.66717
R2229 iovdd.n1309 iovdd.n305 5.66717
R2230 iovdd.n1309 iovdd.n304 5.66717
R2231 iovdd.n1309 iovdd.n302 5.66717
R2232 iovdd.n1309 iovdd.n299 5.66717
R2233 iovdd.n1309 iovdd.n361 5.66717
R2234 iovdd.n1229 iovdd.n567 5.66717
R2235 iovdd.n1229 iovdd.n854 5.66717
R2236 iovdd.n1230 iovdd.n1229 5.66717
R2237 iovdd.n1229 iovdd.n852 5.66717
R2238 iovdd.n1229 iovdd.n848 5.66717
R2239 iovdd.n1229 iovdd.n844 5.66717
R2240 iovdd.n1229 iovdd.n842 5.66717
R2241 iovdd.n1229 iovdd.n840 5.66717
R2242 iovdd.n1229 iovdd.n839 5.66717
R2243 iovdd.n1229 iovdd.n837 5.66717
R2244 iovdd.n1229 iovdd.n835 5.66717
R2245 iovdd.n1229 iovdd.n833 5.66717
R2246 iovdd.n1229 iovdd.n831 5.66717
R2247 iovdd.n1229 iovdd.n830 5.66717
R2248 iovdd.n1229 iovdd.n828 5.66717
R2249 iovdd.n1229 iovdd.n826 5.66717
R2250 iovdd.n1229 iovdd.n824 5.66717
R2251 iovdd.n1229 iovdd.n823 5.66717
R2252 iovdd.n1229 iovdd.n821 5.66717
R2253 iovdd.n1229 iovdd.n819 5.66717
R2254 iovdd.n1229 iovdd.n817 5.66717
R2255 iovdd.n1229 iovdd.n815 5.66717
R2256 iovdd.n1229 iovdd.n814 5.66717
R2257 iovdd.n1229 iovdd.n812 5.66717
R2258 iovdd.n1229 iovdd.n810 5.66717
R2259 iovdd.n1229 iovdd.n808 5.66717
R2260 iovdd.n1229 iovdd.n806 5.66717
R2261 iovdd.n1229 iovdd.n805 5.66717
R2262 iovdd.n1229 iovdd.n803 5.66717
R2263 iovdd.n1229 iovdd.n801 5.66717
R2264 iovdd.n1229 iovdd.n799 5.66717
R2265 iovdd.n1229 iovdd.n797 5.66717
R2266 iovdd.n1229 iovdd.n796 5.66717
R2267 iovdd.n1229 iovdd.n794 5.66717
R2268 iovdd.n1229 iovdd.n792 5.66717
R2269 iovdd.t0 iovdd.n43 5.66717
R2270 iovdd.t0 iovdd.n4 5.66717
R2271 iovdd.t0 iovdd.n42 5.66717
R2272 iovdd.t0 iovdd.n40 5.66717
R2273 iovdd.t0 iovdd.n39 5.66717
R2274 iovdd.t0 iovdd.n37 5.66717
R2275 iovdd.t0 iovdd.n36 5.66717
R2276 iovdd.t0 iovdd.n34 5.66717
R2277 iovdd.t0 iovdd.n33 5.66717
R2278 iovdd.t0 iovdd.n31 5.66717
R2279 iovdd.t0 iovdd.n30 5.66717
R2280 iovdd.t0 iovdd.n28 5.66717
R2281 iovdd.t0 iovdd.n27 5.66717
R2282 iovdd.t0 iovdd.n23 5.66717
R2283 iovdd.t0 iovdd.n22 5.66717
R2284 iovdd.t0 iovdd.n20 5.66717
R2285 iovdd.t0 iovdd.n19 5.66717
R2286 iovdd.t0 iovdd.n17 5.66717
R2287 iovdd.t0 iovdd.n16 5.66717
R2288 iovdd.t0 iovdd.n13 5.66717
R2289 iovdd.t0 iovdd.n12 5.66717
R2290 iovdd.t0 iovdd.n11 5.66717
R2291 iovdd.t0 iovdd.n10 5.66717
R2292 iovdd.t0 iovdd.n9 5.66717
R2293 iovdd.t0 iovdd.n7 5.66717
R2294 iovdd.t0 iovdd.n5 5.66717
R2295 iovdd.n1359 iovdd.n108 5.66717
R2296 iovdd.n1359 iovdd.n106 5.66717
R2297 iovdd.n1359 iovdd.n105 5.66717
R2298 iovdd.n1359 iovdd.n103 5.66717
R2299 iovdd.n1359 iovdd.n101 5.66717
R2300 iovdd.n1359 iovdd.n99 5.66717
R2301 iovdd.n1359 iovdd.n97 5.66717
R2302 iovdd.n1359 iovdd.n96 5.66717
R2303 iovdd.n1359 iovdd.n94 5.66717
R2304 iovdd.n1359 iovdd.n92 5.66717
R2305 iovdd.n1359 iovdd.n90 5.66717
R2306 iovdd.n1359 iovdd.n88 5.66717
R2307 iovdd.n1359 iovdd.n87 5.66717
R2308 iovdd.n1359 iovdd.n85 5.66717
R2309 iovdd.n1359 iovdd.n83 5.66717
R2310 iovdd.n1359 iovdd.n81 5.66717
R2311 iovdd.n1359 iovdd.n80 5.66717
R2312 iovdd.n1359 iovdd.n78 5.66717
R2313 iovdd.n1359 iovdd.n76 5.66717
R2314 iovdd.n1359 iovdd.n74 5.66717
R2315 iovdd.n1359 iovdd.n72 5.66717
R2316 iovdd.n1359 iovdd.n71 5.66717
R2317 iovdd.n1359 iovdd.n69 5.66717
R2318 iovdd.n1359 iovdd.n67 5.66717
R2319 iovdd.n1359 iovdd.n65 5.66717
R2320 iovdd.n1359 iovdd.n63 5.66717
R2321 iovdd.n1359 iovdd.n62 5.66717
R2322 iovdd.n1359 iovdd.n60 5.66717
R2323 iovdd.n1359 iovdd.n58 5.66717
R2324 iovdd.n1359 iovdd.n56 5.66717
R2325 iovdd.n1359 iovdd.n54 5.66717
R2326 iovdd.n1359 iovdd.n53 5.66717
R2327 iovdd.n1359 iovdd.n51 5.66717
R2328 iovdd.n1359 iovdd.n46 5.66717
R2329 iovdd.n1359 iovdd.n110 5.66717
R2330 iovdd.n1359 iovdd.n45 5.66717
R2331 iovdd.n1359 iovdd.n1358 5.66717
R2332 iovdd.n289 iovdd.n288 5.66717
R2333 iovdd.n288 iovdd.n277 5.66717
R2334 iovdd.n1310 iovdd.n1309 5.66717
R2335 iovdd.n3 iovdd.n0 5.66717
R2336 iovdd.n861 iovdd.n3 5.66717
R2337 iovdd.n1229 iovdd.n1228 5.66717
R2338 iovdd.n550 iovdd.n548 4.50058
R2339 iovdd.n297 iovdd.n248 4.50058
R2340 iovdd.n1222 iovdd.n1089 4.50058
R2341 iovdd.n1226 iovdd.n864 4.50058
R2342 iovdd.n1329 iovdd.n113 4.50058
R2343 iovdd.n1297 iovdd.n1296 4.50058
R2344 iovdd.n781 iovdd.n387 4.50058
R2345 iovdd.n547 iovdd.n480 4.49246
R2346 iovdd.n477 iovdd.n431 4.49246
R2347 iovdd.n1313 iovdd.n271 4.49246
R2348 iovdd.n481 iovdd.n431 4.49246
R2349 iovdd.n1313 iovdd.n270 4.49246
R2350 iovdd.n484 iovdd.n431 4.49246
R2351 iovdd.n1313 iovdd.n269 4.49246
R2352 iovdd.n487 iovdd.n431 4.49246
R2353 iovdd.n1313 iovdd.n268 4.49246
R2354 iovdd.n490 iovdd.n431 4.49246
R2355 iovdd.n1313 iovdd.n267 4.49246
R2356 iovdd.n493 iovdd.n431 4.49246
R2357 iovdd.n1313 iovdd.n266 4.49246
R2358 iovdd.n496 iovdd.n431 4.49246
R2359 iovdd.n1313 iovdd.n265 4.49246
R2360 iovdd.n499 iovdd.n431 4.49246
R2361 iovdd.n1313 iovdd.n264 4.49246
R2362 iovdd.n502 iovdd.n431 4.49246
R2363 iovdd.n1313 iovdd.n263 4.49246
R2364 iovdd.n505 iovdd.n431 4.49246
R2365 iovdd.n1313 iovdd.n262 4.49246
R2366 iovdd.n508 iovdd.n431 4.49246
R2367 iovdd.n1313 iovdd.n261 4.49246
R2368 iovdd.n511 iovdd.n431 4.49246
R2369 iovdd.n1313 iovdd.n260 4.49246
R2370 iovdd.n514 iovdd.n431 4.49246
R2371 iovdd.n1313 iovdd.n259 4.49246
R2372 iovdd.n517 iovdd.n431 4.49246
R2373 iovdd.n1313 iovdd.n258 4.49246
R2374 iovdd.n520 iovdd.n431 4.49246
R2375 iovdd.n1313 iovdd.n257 4.49246
R2376 iovdd.n523 iovdd.n431 4.49246
R2377 iovdd.n1313 iovdd.n256 4.49246
R2378 iovdd.n526 iovdd.n431 4.49246
R2379 iovdd.n1313 iovdd.n255 4.49246
R2380 iovdd.n529 iovdd.n431 4.49246
R2381 iovdd.n1313 iovdd.n254 4.49246
R2382 iovdd.n532 iovdd.n431 4.49246
R2383 iovdd.n1313 iovdd.n253 4.49246
R2384 iovdd.n535 iovdd.n431 4.49246
R2385 iovdd.n1313 iovdd.n252 4.49246
R2386 iovdd.n538 iovdd.n431 4.49246
R2387 iovdd.n1313 iovdd.n251 4.49246
R2388 iovdd.n541 iovdd.n431 4.49246
R2389 iovdd.n1313 iovdd.n250 4.49246
R2390 iovdd.n544 iovdd.n431 4.49246
R2391 iovdd.n1313 iovdd.n249 4.49246
R2392 iovdd.n431 iovdd.n274 4.49246
R2393 iovdd.n547 iovdd.n276 4.49246
R2394 iovdd.n1218 iovdd.n1217 4.49246
R2395 iovdd.n1223 iovdd.n1087 4.49246
R2396 iovdd.n1218 iovdd.n1216 4.49246
R2397 iovdd.n1223 iovdd.n1086 4.49246
R2398 iovdd.n1218 iovdd.n1215 4.49246
R2399 iovdd.n1223 iovdd.n1085 4.49246
R2400 iovdd.n1218 iovdd.n1214 4.49246
R2401 iovdd.n1223 iovdd.n1084 4.49246
R2402 iovdd.n1218 iovdd.n1213 4.49246
R2403 iovdd.n1223 iovdd.n1083 4.49246
R2404 iovdd.n1218 iovdd.n1212 4.49246
R2405 iovdd.n1223 iovdd.n1082 4.49246
R2406 iovdd.n1218 iovdd.n1211 4.49246
R2407 iovdd.n1223 iovdd.n1081 4.49246
R2408 iovdd.n1218 iovdd.n1210 4.49246
R2409 iovdd.n1223 iovdd.n1080 4.49246
R2410 iovdd.n1218 iovdd.n1209 4.49246
R2411 iovdd.n1223 iovdd.n1079 4.49246
R2412 iovdd.n1218 iovdd.n1208 4.49246
R2413 iovdd.n1223 iovdd.n1078 4.49246
R2414 iovdd.n1218 iovdd.n1207 4.49246
R2415 iovdd.n1223 iovdd.n1077 4.49246
R2416 iovdd.n1218 iovdd.n1206 4.49246
R2417 iovdd.n1223 iovdd.n1076 4.49246
R2418 iovdd.n1218 iovdd.n1205 4.49246
R2419 iovdd.n1223 iovdd.n1075 4.49246
R2420 iovdd.n1218 iovdd.n1204 4.49246
R2421 iovdd.n1223 iovdd.n1074 4.49246
R2422 iovdd.n1218 iovdd.n1203 4.49246
R2423 iovdd.n1223 iovdd.n1073 4.49246
R2424 iovdd.n1218 iovdd.n1202 4.49246
R2425 iovdd.n1223 iovdd.n1072 4.49246
R2426 iovdd.n1218 iovdd.n1201 4.49246
R2427 iovdd.n1223 iovdd.n1071 4.49246
R2428 iovdd.n1218 iovdd.n1200 4.49246
R2429 iovdd.n1223 iovdd.n1070 4.49246
R2430 iovdd.n1218 iovdd.n1199 4.49246
R2431 iovdd.n1223 iovdd.n1069 4.49246
R2432 iovdd.n1218 iovdd.n1198 4.49246
R2433 iovdd.n1223 iovdd.n1068 4.49246
R2434 iovdd.n1218 iovdd.n1197 4.49246
R2435 iovdd.n1223 iovdd.n1067 4.49246
R2436 iovdd.n1218 iovdd.n1196 4.49246
R2437 iovdd.n1223 iovdd.n1066 4.49246
R2438 iovdd.n1218 iovdd.n1195 4.49246
R2439 iovdd.n1223 iovdd.n1065 4.49246
R2440 iovdd.n1224 iovdd.n1223 4.49246
R2441 iovdd.n117 iovdd.n116 4.49246
R2442 iovdd.n1353 iovdd.n114 4.49246
R2443 iovdd.n166 iovdd.n115 4.49246
R2444 iovdd.n1353 iovdd.n1330 4.49246
R2445 iovdd.n169 iovdd.n115 4.49246
R2446 iovdd.n1353 iovdd.n1331 4.49246
R2447 iovdd.n172 iovdd.n115 4.49246
R2448 iovdd.n1353 iovdd.n1332 4.49246
R2449 iovdd.n175 iovdd.n115 4.49246
R2450 iovdd.n1353 iovdd.n1333 4.49246
R2451 iovdd.n178 iovdd.n115 4.49246
R2452 iovdd.n1353 iovdd.n1334 4.49246
R2453 iovdd.n181 iovdd.n115 4.49246
R2454 iovdd.n1353 iovdd.n1335 4.49246
R2455 iovdd.n184 iovdd.n115 4.49246
R2456 iovdd.n1353 iovdd.n1336 4.49246
R2457 iovdd.n187 iovdd.n115 4.49246
R2458 iovdd.n1353 iovdd.n1337 4.49246
R2459 iovdd.n190 iovdd.n115 4.49246
R2460 iovdd.n1353 iovdd.n1338 4.49246
R2461 iovdd.n193 iovdd.n115 4.49246
R2462 iovdd.n1353 iovdd.n1339 4.49246
R2463 iovdd.n196 iovdd.n115 4.49246
R2464 iovdd.n1353 iovdd.n1340 4.49246
R2465 iovdd.n199 iovdd.n115 4.49246
R2466 iovdd.n1353 iovdd.n1341 4.49246
R2467 iovdd.n202 iovdd.n115 4.49246
R2468 iovdd.n1353 iovdd.n1342 4.49246
R2469 iovdd.n205 iovdd.n115 4.49246
R2470 iovdd.n1353 iovdd.n1343 4.49246
R2471 iovdd.n208 iovdd.n115 4.49246
R2472 iovdd.n1353 iovdd.n1344 4.49246
R2473 iovdd.n211 iovdd.n115 4.49246
R2474 iovdd.n1353 iovdd.n1345 4.49246
R2475 iovdd.n214 iovdd.n115 4.49246
R2476 iovdd.n1353 iovdd.n1346 4.49246
R2477 iovdd.n217 iovdd.n115 4.49246
R2478 iovdd.n1353 iovdd.n1347 4.49246
R2479 iovdd.n220 iovdd.n115 4.49246
R2480 iovdd.n1353 iovdd.n1348 4.49246
R2481 iovdd.n223 iovdd.n115 4.49246
R2482 iovdd.n1353 iovdd.n1349 4.49246
R2483 iovdd.n226 iovdd.n115 4.49246
R2484 iovdd.n1353 iovdd.n1350 4.49246
R2485 iovdd.n229 iovdd.n115 4.49246
R2486 iovdd.n1353 iovdd.n1351 4.49246
R2487 iovdd.n232 iovdd.n115 4.49246
R2488 iovdd.n1353 iovdd.n1352 4.49246
R2489 iovdd.n237 iovdd.n115 4.49246
R2490 iovdd.n1304 iovdd.n401 4.49246
R2491 iovdd.n1298 iovdd.n389 4.49246
R2492 iovdd.n1301 iovdd.n1281 4.49246
R2493 iovdd.n402 iovdd.n389 4.49246
R2494 iovdd.n1301 iovdd.n1280 4.49246
R2495 iovdd.n405 iovdd.n389 4.49246
R2496 iovdd.n1301 iovdd.n1279 4.49246
R2497 iovdd.n408 iovdd.n389 4.49246
R2498 iovdd.n1302 iovdd.n1301 4.49246
R2499 iovdd.n411 iovdd.n389 4.49246
R2500 iovdd.n1301 iovdd.n390 4.49246
R2501 iovdd.n1249 iovdd.n559 4.49246
R2502 iovdd.n1264 iovdd.n560 4.49246
R2503 iovdd.n1252 iovdd.n559 4.49246
R2504 iovdd.n1264 iovdd.n561 4.49246
R2505 iovdd.n1255 iovdd.n559 4.49246
R2506 iovdd.n1264 iovdd.n562 4.49246
R2507 iovdd.n1258 iovdd.n559 4.49246
R2508 iovdd.n1264 iovdd.n563 4.49246
R2509 iovdd.n566 iovdd.n559 4.49246
R2510 iovdd.n1264 iovdd.n1263 4.49246
R2511 iovdd.n564 iovdd.n559 4.49246
R2512 iovdd.n785 iovdd.n774 4.49246
R2513 iovdd.n1236 iovdd.n775 4.49246
R2514 iovdd.n787 iovdd.n774 4.49246
R2515 iovdd.n1236 iovdd.n776 4.49246
R2516 iovdd.n789 iovdd.n774 4.49246
R2517 iovdd.n1236 iovdd.n777 4.49246
R2518 iovdd.n779 iovdd.n774 4.49246
R2519 iovdd.n1236 iovdd.n1235 4.49246
R2520 iovdd.n774 iovdd.n569 4.49246
R2521 iovdd.n1233 iovdd.n568 4.49246
R2522 iovdd.n1236 iovdd.n770 4.49246
R2523 iovdd.n298 iovdd.n272 3.0005
R2524 iovdd.n1262 iovdd.n1240 3.0005
R2525 iovdd.n483 iovdd.n482 3.0005
R2526 iovdd.n474 iovdd.n473 3.0005
R2527 iovdd.n472 iovdd.n471 3.0005
R2528 iovdd.n470 iovdd.n469 3.0005
R2529 iovdd.n468 iovdd.n467 3.0005
R2530 iovdd.n498 iovdd.n497 3.0005
R2531 iovdd.n501 iovdd.n500 3.0005
R2532 iovdd.n504 iovdd.n503 3.0005
R2533 iovdd.n507 iovdd.n506 3.0005
R2534 iovdd.n510 iovdd.n509 3.0005
R2535 iovdd.n458 iovdd.n457 3.0005
R2536 iovdd.n456 iovdd.n455 3.0005
R2537 iovdd.n454 iovdd.n453 3.0005
R2538 iovdd.n452 iovdd.n451 3.0005
R2539 iovdd.n450 iovdd.n449 3.0005
R2540 iovdd.n525 iovdd.n524 3.0005
R2541 iovdd.n528 iovdd.n527 3.0005
R2542 iovdd.n531 iovdd.n530 3.0005
R2543 iovdd.n534 iovdd.n533 3.0005
R2544 iovdd.n440 iovdd.n439 3.0005
R2545 iovdd.n438 iovdd.n437 3.0005
R2546 iovdd.n436 iovdd.n435 3.0005
R2547 iovdd.n434 iovdd.n433 3.0005
R2548 iovdd.n550 iovdd.n549 3.0005
R2549 iovdd.n430 iovdd.n429 3.0005
R2550 iovdd.n556 iovdd.n427 3.0005
R2551 iovdd.n424 iovdd.n423 3.0005
R2552 iovdd.n1248 iovdd.n1247 3.0005
R2553 iovdd.n1254 iovdd.n1253 3.0005
R2554 iovdd.n1257 iovdd.n1256 3.0005
R2555 iovdd.n1260 iovdd.n1259 3.0005
R2556 iovdd.n1242 iovdd.n1241 3.0005
R2557 iovdd.n1244 iovdd.n1243 3.0005
R2558 iovdd.n1246 iovdd.n1245 3.0005
R2559 iovdd.n1251 iovdd.n1250 3.0005
R2560 iovdd.n557 iovdd.n426 3.0005
R2561 iovdd.n555 iovdd.n428 3.0005
R2562 iovdd.n551 iovdd.n432 3.0005
R2563 iovdd.n546 iovdd.n545 3.0005
R2564 iovdd.n543 iovdd.n542 3.0005
R2565 iovdd.n540 iovdd.n539 3.0005
R2566 iovdd.n537 iovdd.n536 3.0005
R2567 iovdd.n442 iovdd.n441 3.0005
R2568 iovdd.n444 iovdd.n443 3.0005
R2569 iovdd.n446 iovdd.n445 3.0005
R2570 iovdd.n448 iovdd.n447 3.0005
R2571 iovdd.n522 iovdd.n521 3.0005
R2572 iovdd.n519 iovdd.n518 3.0005
R2573 iovdd.n516 iovdd.n515 3.0005
R2574 iovdd.n513 iovdd.n512 3.0005
R2575 iovdd.n460 iovdd.n459 3.0005
R2576 iovdd.n462 iovdd.n461 3.0005
R2577 iovdd.n464 iovdd.n463 3.0005
R2578 iovdd.n466 iovdd.n465 3.0005
R2579 iovdd.n495 iovdd.n494 3.0005
R2580 iovdd.n492 iovdd.n491 3.0005
R2581 iovdd.n489 iovdd.n488 3.0005
R2582 iovdd.n486 iovdd.n485 3.0005
R2583 iovdd.n476 iovdd.n475 3.0005
R2584 iovdd.n479 iovdd.n478 3.0005
R2585 iovdd.n300 iovdd.n273 3.0005
R2586 iovdd.n552 iovdd.n551 3.0005
R2587 iovdd.n553 iovdd.n430 3.0005
R2588 iovdd.n555 iovdd.n554 3.0005
R2589 iovdd.n556 iovdd.n425 3.0005
R2590 iovdd.n558 iovdd.n557 3.0005
R2591 iovdd.n1194 iovdd.n1090 3.0005
R2592 iovdd.n1192 iovdd.n1190 3.0005
R2593 iovdd.n1189 iovdd.n1182 3.0005
R2594 iovdd.n1188 iovdd.n1187 3.0005
R2595 iovdd.n1185 iovdd.n1183 3.0005
R2596 iovdd.n1306 iovdd.n387 3.0005
R2597 iovdd.n1306 iovdd.n388 3.0005
R2598 iovdd.n772 iovdd.n565 3.0005
R2599 iovdd.n773 iovdd.n772 3.0005
R2600 iovdd.n862 iovdd.n859 3.0005
R2601 iovdd.n1238 iovdd.n1237 3.0005
R2602 iovdd.n855 iovdd.n778 3.0005
R2603 iovdd.n1234 iovdd.n780 3.0005
R2604 iovdd.n853 iovdd.n782 3.0005
R2605 iovdd.n1232 iovdd.n1231 3.0005
R2606 iovdd.n791 iovdd.n783 3.0005
R2607 iovdd.n851 iovdd.n788 3.0005
R2608 iovdd.n849 iovdd.n784 3.0005
R2609 iovdd.n847 iovdd.n786 3.0005
R2610 iovdd.n845 iovdd.n771 3.0005
R2611 iovdd.n1185 iovdd.n1184 3.0005
R2612 iovdd.n1187 iovdd.n1186 3.0005
R2613 iovdd.n1182 iovdd.n1181 3.0005
R2614 iovdd.n1192 iovdd.n1191 3.0005
R2615 iovdd.n1194 iovdd.n1193 3.0005
R2616 iovdd.n1220 iovdd.n1219 3.0005
R2617 iovdd.n1092 iovdd.n1091 3.0005
R2618 iovdd.n1180 iovdd.n1179 3.0005
R2619 iovdd.n1094 iovdd.n1093 3.0005
R2620 iovdd.n1178 iovdd.n1177 3.0005
R2621 iovdd.n1096 iovdd.n1095 3.0005
R2622 iovdd.n1176 iovdd.n1175 3.0005
R2623 iovdd.n1098 iovdd.n1097 3.0005
R2624 iovdd.n1174 iovdd.n1173 3.0005
R2625 iovdd.n1100 iovdd.n1099 3.0005
R2626 iovdd.n1172 iovdd.n1171 3.0005
R2627 iovdd.n1102 iovdd.n1101 3.0005
R2628 iovdd.n1170 iovdd.n1169 3.0005
R2629 iovdd.n1104 iovdd.n1103 3.0005
R2630 iovdd.n1168 iovdd.n1167 3.0005
R2631 iovdd.n1106 iovdd.n1105 3.0005
R2632 iovdd.n1166 iovdd.n1165 3.0005
R2633 iovdd.n1108 iovdd.n1107 3.0005
R2634 iovdd.n1164 iovdd.n1163 3.0005
R2635 iovdd.n1110 iovdd.n1109 3.0005
R2636 iovdd.n1162 iovdd.n1161 3.0005
R2637 iovdd.n1112 iovdd.n1111 3.0005
R2638 iovdd.n1160 iovdd.n1159 3.0005
R2639 iovdd.n1114 iovdd.n1113 3.0005
R2640 iovdd.n1158 iovdd.n1157 3.0005
R2641 iovdd.n1116 iovdd.n1115 3.0005
R2642 iovdd.n1156 iovdd.n1155 3.0005
R2643 iovdd.n1118 iovdd.n1117 3.0005
R2644 iovdd.n1154 iovdd.n1153 3.0005
R2645 iovdd.n1120 iovdd.n1119 3.0005
R2646 iovdd.n1152 iovdd.n1151 3.0005
R2647 iovdd.n1122 iovdd.n1121 3.0005
R2648 iovdd.n1150 iovdd.n1149 3.0005
R2649 iovdd.n1124 iovdd.n1123 3.0005
R2650 iovdd.n1148 iovdd.n1147 3.0005
R2651 iovdd.n1126 iovdd.n1125 3.0005
R2652 iovdd.n1146 iovdd.n1145 3.0005
R2653 iovdd.n1128 iovdd.n1127 3.0005
R2654 iovdd.n1144 iovdd.n1143 3.0005
R2655 iovdd.n1130 iovdd.n1129 3.0005
R2656 iovdd.n1142 iovdd.n1141 3.0005
R2657 iovdd.n1132 iovdd.n1131 3.0005
R2658 iovdd.n1140 iovdd.n1139 3.0005
R2659 iovdd.n1134 iovdd.n1133 3.0005
R2660 iovdd.n1138 iovdd.n1137 3.0005
R2661 iovdd.n1136 iovdd.n1135 3.0005
R2662 iovdd.n1089 iovdd.n1088 3.0005
R2663 iovdd.n165 iovdd.n112 3.0005
R2664 iovdd.n396 iovdd.n395 3.0005
R2665 iovdd.n407 iovdd.n406 3.0005
R2666 iovdd.n398 iovdd.n397 3.0005
R2667 iovdd.n404 iovdd.n403 3.0005
R2668 iovdd.n400 iovdd.n399 3.0005
R2669 iovdd.n1300 iovdd.n1299 3.0005
R2670 iovdd.n1296 iovdd.n1282 3.0005
R2671 iovdd.n1295 iovdd.n1283 3.0005
R2672 iovdd.n1285 iovdd.n1284 3.0005
R2673 iovdd.n1291 iovdd.n1288 3.0005
R2674 iovdd.n1290 iovdd.n1289 3.0005
R2675 iovdd.n236 iovdd.n235 3.0005
R2676 iovdd.n1354 iovdd.n238 3.0005
R2677 iovdd.n120 iovdd.n119 3.0005
R2678 iovdd.n234 iovdd.n233 3.0005
R2679 iovdd.n122 iovdd.n121 3.0005
R2680 iovdd.n231 iovdd.n230 3.0005
R2681 iovdd.n124 iovdd.n123 3.0005
R2682 iovdd.n228 iovdd.n227 3.0005
R2683 iovdd.n126 iovdd.n125 3.0005
R2684 iovdd.n225 iovdd.n224 3.0005
R2685 iovdd.n128 iovdd.n127 3.0005
R2686 iovdd.n222 iovdd.n221 3.0005
R2687 iovdd.n130 iovdd.n129 3.0005
R2688 iovdd.n219 iovdd.n218 3.0005
R2689 iovdd.n132 iovdd.n131 3.0005
R2690 iovdd.n216 iovdd.n215 3.0005
R2691 iovdd.n134 iovdd.n133 3.0005
R2692 iovdd.n213 iovdd.n212 3.0005
R2693 iovdd.n136 iovdd.n135 3.0005
R2694 iovdd.n210 iovdd.n209 3.0005
R2695 iovdd.n138 iovdd.n137 3.0005
R2696 iovdd.n207 iovdd.n206 3.0005
R2697 iovdd.n140 iovdd.n139 3.0005
R2698 iovdd.n204 iovdd.n203 3.0005
R2699 iovdd.n142 iovdd.n141 3.0005
R2700 iovdd.n201 iovdd.n200 3.0005
R2701 iovdd.n144 iovdd.n143 3.0005
R2702 iovdd.n198 iovdd.n197 3.0005
R2703 iovdd.n146 iovdd.n145 3.0005
R2704 iovdd.n195 iovdd.n194 3.0005
R2705 iovdd.n148 iovdd.n147 3.0005
R2706 iovdd.n192 iovdd.n191 3.0005
R2707 iovdd.n150 iovdd.n149 3.0005
R2708 iovdd.n189 iovdd.n188 3.0005
R2709 iovdd.n152 iovdd.n151 3.0005
R2710 iovdd.n186 iovdd.n185 3.0005
R2711 iovdd.n154 iovdd.n153 3.0005
R2712 iovdd.n183 iovdd.n182 3.0005
R2713 iovdd.n156 iovdd.n155 3.0005
R2714 iovdd.n180 iovdd.n179 3.0005
R2715 iovdd.n158 iovdd.n157 3.0005
R2716 iovdd.n177 iovdd.n176 3.0005
R2717 iovdd.n160 iovdd.n159 3.0005
R2718 iovdd.n174 iovdd.n173 3.0005
R2719 iovdd.n162 iovdd.n161 3.0005
R2720 iovdd.n171 iovdd.n170 3.0005
R2721 iovdd.n164 iovdd.n163 3.0005
R2722 iovdd.n168 iovdd.n167 3.0005
R2723 iovdd.n1303 iovdd.n412 3.0005
R2724 iovdd.n1306 iovdd.n1305 3.0005
R2725 iovdd.n772 iovdd.n392 3.0005
R2726 iovdd.n394 iovdd.n393 3.0005
R2727 iovdd.n410 iovdd.n409 3.0005
R2728 iovdd.n1286 iovdd.n236 3.0005
R2729 iovdd.n1290 iovdd.n1287 3.0005
R2730 iovdd.n1292 iovdd.n1291 3.0005
R2731 iovdd.n1293 iovdd.n1285 3.0005
R2732 iovdd.n1295 iovdd.n1294 3.0005
R2733 iovdd.t0 iovdd.n24 2.83433
R2734 iovdd.t0 iovdd.n21 2.83433
R2735 iovdd.t0 iovdd.n18 2.83433
R2736 iovdd.t0 iovdd.n15 2.83433
R2737 iovdd.t0 iovdd.n2 2.83433
R2738 iovdd.n1361 iovdd.t0 2.83433
R2739 iovdd.t0 iovdd.n6 2.83433
R2740 iovdd.t0 iovdd.n41 2.83433
R2741 iovdd.t0 iovdd.n38 2.83433
R2742 iovdd.t0 iovdd.n35 2.83433
R2743 iovdd.t0 iovdd.n32 2.83433
R2744 iovdd.t0 iovdd.n29 2.83433
R2745 iovdd.t0 iovdd.n26 2.83433
R2746 iovdd.n1309 iovdd.n360 2.82693
R2747 iovdd.n1309 iovdd.n358 2.82693
R2748 iovdd.n1309 iovdd.n355 2.82693
R2749 iovdd.n1309 iovdd.n353 2.82693
R2750 iovdd.n1309 iovdd.n351 2.82693
R2751 iovdd.n1309 iovdd.n349 2.82693
R2752 iovdd.n1309 iovdd.n346 2.82693
R2753 iovdd.n1309 iovdd.n344 2.82693
R2754 iovdd.n1309 iovdd.n342 2.82693
R2755 iovdd.n1309 iovdd.n340 2.82693
R2756 iovdd.n1309 iovdd.n337 2.82693
R2757 iovdd.n1309 iovdd.n335 2.82693
R2758 iovdd.n1309 iovdd.n333 2.82693
R2759 iovdd.n1309 iovdd.n331 2.82693
R2760 iovdd.n1309 iovdd.n328 2.82693
R2761 iovdd.n1309 iovdd.n326 2.82693
R2762 iovdd.n1309 iovdd.n324 2.82693
R2763 iovdd.n1309 iovdd.n321 2.82693
R2764 iovdd.n1309 iovdd.n319 2.82693
R2765 iovdd.n1309 iovdd.n317 2.82693
R2766 iovdd.n1309 iovdd.n315 2.82693
R2767 iovdd.n1309 iovdd.n312 2.82693
R2768 iovdd.n1309 iovdd.n310 2.82693
R2769 iovdd.n1309 iovdd.n308 2.82693
R2770 iovdd.n1309 iovdd.n306 2.82693
R2771 iovdd.n1309 iovdd.n303 2.82693
R2772 iovdd.n1309 iovdd.n301 2.82693
R2773 iovdd.n1229 iovdd.n856 2.82693
R2774 iovdd.n1229 iovdd.n790 2.82693
R2775 iovdd.n1229 iovdd.n850 2.82693
R2776 iovdd.n1229 iovdd.n846 2.82693
R2777 iovdd.n1229 iovdd.n843 2.82693
R2778 iovdd.n1229 iovdd.n841 2.82693
R2779 iovdd.n1229 iovdd.n838 2.82693
R2780 iovdd.n1229 iovdd.n836 2.82693
R2781 iovdd.n1229 iovdd.n834 2.82693
R2782 iovdd.n1229 iovdd.n832 2.82693
R2783 iovdd.n1229 iovdd.n829 2.82693
R2784 iovdd.n1229 iovdd.n827 2.82693
R2785 iovdd.n1229 iovdd.n825 2.82693
R2786 iovdd.n1229 iovdd.n822 2.82693
R2787 iovdd.n1229 iovdd.n820 2.82693
R2788 iovdd.n1229 iovdd.n818 2.82693
R2789 iovdd.n1229 iovdd.n816 2.82693
R2790 iovdd.n1229 iovdd.n813 2.82693
R2791 iovdd.n1229 iovdd.n811 2.82693
R2792 iovdd.n1229 iovdd.n809 2.82693
R2793 iovdd.n1229 iovdd.n807 2.82693
R2794 iovdd.n1229 iovdd.n804 2.82693
R2795 iovdd.n1229 iovdd.n802 2.82693
R2796 iovdd.n1229 iovdd.n800 2.82693
R2797 iovdd.n1229 iovdd.n798 2.82693
R2798 iovdd.n1229 iovdd.n795 2.82693
R2799 iovdd.n1229 iovdd.n793 2.82693
R2800 iovdd.n1359 iovdd.n109 2.82693
R2801 iovdd.n1359 iovdd.n107 2.82693
R2802 iovdd.n1359 iovdd.n104 2.82693
R2803 iovdd.n1359 iovdd.n102 2.82693
R2804 iovdd.n1359 iovdd.n100 2.82693
R2805 iovdd.n1359 iovdd.n98 2.82693
R2806 iovdd.n1359 iovdd.n95 2.82693
R2807 iovdd.n1359 iovdd.n93 2.82693
R2808 iovdd.n1359 iovdd.n91 2.82693
R2809 iovdd.n1359 iovdd.n89 2.82693
R2810 iovdd.n1359 iovdd.n86 2.82693
R2811 iovdd.n1359 iovdd.n84 2.82693
R2812 iovdd.n1359 iovdd.n82 2.82693
R2813 iovdd.n1359 iovdd.n79 2.82693
R2814 iovdd.n1359 iovdd.n77 2.82693
R2815 iovdd.n1359 iovdd.n75 2.82693
R2816 iovdd.n1359 iovdd.n73 2.82693
R2817 iovdd.n1359 iovdd.n70 2.82693
R2818 iovdd.n1359 iovdd.n68 2.82693
R2819 iovdd.n1359 iovdd.n66 2.82693
R2820 iovdd.n1359 iovdd.n64 2.82693
R2821 iovdd.n1359 iovdd.n61 2.82693
R2822 iovdd.n1359 iovdd.n59 2.82693
R2823 iovdd.n1359 iovdd.n57 2.82693
R2824 iovdd.n1359 iovdd.n55 2.82693
R2825 iovdd.n1359 iovdd.n52 2.82693
R2826 iovdd.n1359 iovdd.n50 2.82693
R2827 iovdd.n279 iovdd.n278 2.82693
R2828 iovdd.n281 iovdd.n280 2.82693
R2829 iovdd.n283 iovdd.n282 2.82693
R2830 iovdd.n285 iovdd.n284 2.82693
R2831 iovdd.n287 iovdd.n286 2.82693
R2832 iovdd.n296 iovdd.n291 2.82693
R2833 iovdd.n295 iovdd.n292 2.82693
R2834 iovdd.n294 iovdd.n293 2.82693
R2835 iovdd.n14 iovdd.n1 2.82693
R2836 iovdd.n1363 iovdd.n1362 2.82693
R2837 iovdd.n944 iovdd.n937 0.826084
R2838 iovdd.n649 iovdd.n642 0.826084
R2839 iovdd.n1326 iovdd.n1325 0.822133
R2840 iovdd.n1275 iovdd.n415 0.822133
R2841 iovdd.n943 iovdd.n942 0.818682
R2842 iovdd.n938 iovdd.n936 0.818682
R2843 iovdd.n948 iovdd.n947 0.818682
R2844 iovdd.n949 iovdd.n929 0.818682
R2845 iovdd.n958 iovdd.n957 0.818682
R2846 iovdd.n931 iovdd.n927 0.818682
R2847 iovdd.n963 iovdd.n962 0.818682
R2848 iovdd.n964 iovdd.n920 0.818682
R2849 iovdd.n973 iovdd.n972 0.818682
R2850 iovdd.n922 iovdd.n918 0.818682
R2851 iovdd.n978 iovdd.n977 0.818682
R2852 iovdd.n979 iovdd.n911 0.818682
R2853 iovdd.n988 iovdd.n987 0.818682
R2854 iovdd.n913 iovdd.n909 0.818682
R2855 iovdd.n993 iovdd.n992 0.818682
R2856 iovdd.n994 iovdd.n902 0.818682
R2857 iovdd.n1003 iovdd.n1002 0.818682
R2858 iovdd.n904 iovdd.n900 0.818682
R2859 iovdd.n1008 iovdd.n1007 0.818682
R2860 iovdd.n1009 iovdd.n893 0.818682
R2861 iovdd.n1018 iovdd.n1017 0.818682
R2862 iovdd.n895 iovdd.n891 0.818682
R2863 iovdd.n1023 iovdd.n1022 0.818682
R2864 iovdd.n1024 iovdd.n884 0.818682
R2865 iovdd.n1033 iovdd.n1032 0.818682
R2866 iovdd.n886 iovdd.n882 0.818682
R2867 iovdd.n1038 iovdd.n1037 0.818682
R2868 iovdd.n1039 iovdd.n875 0.818682
R2869 iovdd.n1048 iovdd.n1047 0.818682
R2870 iovdd.n877 iovdd.n873 0.818682
R2871 iovdd.n1053 iovdd.n1052 0.818682
R2872 iovdd.n1054 iovdd.n866 0.818682
R2873 iovdd.n1063 iovdd.n1062 0.818682
R2874 iovdd.n868 iovdd.n246 0.818682
R2875 iovdd.n1316 iovdd.n1315 0.818682
R2876 iovdd.n1318 iovdd.n240 0.818682
R2877 iovdd.n1327 iovdd.n241 0.818682
R2878 iovdd.n1326 iovdd.n118 0.818682
R2879 iovdd.n1328 iovdd.n1327 0.818682
R2880 iovdd.n240 iovdd.n239 0.818682
R2881 iovdd.n1315 iovdd.n1314 0.818682
R2882 iovdd.n247 iovdd.n246 0.818682
R2883 iovdd.n1064 iovdd.n1063 0.818682
R2884 iovdd.n866 iovdd.n865 0.818682
R2885 iovdd.n1052 iovdd.n1051 0.818682
R2886 iovdd.n1050 iovdd.n873 0.818682
R2887 iovdd.n1049 iovdd.n1048 0.818682
R2888 iovdd.n875 iovdd.n874 0.818682
R2889 iovdd.n1037 iovdd.n1036 0.818682
R2890 iovdd.n1035 iovdd.n882 0.818682
R2891 iovdd.n1034 iovdd.n1033 0.818682
R2892 iovdd.n884 iovdd.n883 0.818682
R2893 iovdd.n1022 iovdd.n1021 0.818682
R2894 iovdd.n1020 iovdd.n891 0.818682
R2895 iovdd.n1019 iovdd.n1018 0.818682
R2896 iovdd.n893 iovdd.n892 0.818682
R2897 iovdd.n1007 iovdd.n1006 0.818682
R2898 iovdd.n1005 iovdd.n900 0.818682
R2899 iovdd.n1004 iovdd.n1003 0.818682
R2900 iovdd.n902 iovdd.n901 0.818682
R2901 iovdd.n992 iovdd.n991 0.818682
R2902 iovdd.n990 iovdd.n909 0.818682
R2903 iovdd.n989 iovdd.n988 0.818682
R2904 iovdd.n911 iovdd.n910 0.818682
R2905 iovdd.n977 iovdd.n976 0.818682
R2906 iovdd.n975 iovdd.n918 0.818682
R2907 iovdd.n974 iovdd.n973 0.818682
R2908 iovdd.n920 iovdd.n919 0.818682
R2909 iovdd.n962 iovdd.n961 0.818682
R2910 iovdd.n960 iovdd.n927 0.818682
R2911 iovdd.n959 iovdd.n958 0.818682
R2912 iovdd.n929 iovdd.n928 0.818682
R2913 iovdd.n947 iovdd.n946 0.818682
R2914 iovdd.n945 iovdd.n936 0.818682
R2915 iovdd.n415 iovdd.n391 0.818682
R2916 iovdd.n769 iovdd.n768 0.818682
R2917 iovdd.n571 iovdd.n570 0.818682
R2918 iovdd.n757 iovdd.n756 0.818682
R2919 iovdd.n755 iovdd.n578 0.818682
R2920 iovdd.n754 iovdd.n753 0.818682
R2921 iovdd.n580 iovdd.n579 0.818682
R2922 iovdd.n742 iovdd.n741 0.818682
R2923 iovdd.n740 iovdd.n587 0.818682
R2924 iovdd.n739 iovdd.n738 0.818682
R2925 iovdd.n589 iovdd.n588 0.818682
R2926 iovdd.n727 iovdd.n726 0.818682
R2927 iovdd.n725 iovdd.n596 0.818682
R2928 iovdd.n724 iovdd.n723 0.818682
R2929 iovdd.n598 iovdd.n597 0.818682
R2930 iovdd.n712 iovdd.n711 0.818682
R2931 iovdd.n710 iovdd.n605 0.818682
R2932 iovdd.n709 iovdd.n708 0.818682
R2933 iovdd.n607 iovdd.n606 0.818682
R2934 iovdd.n697 iovdd.n696 0.818682
R2935 iovdd.n695 iovdd.n614 0.818682
R2936 iovdd.n694 iovdd.n693 0.818682
R2937 iovdd.n616 iovdd.n615 0.818682
R2938 iovdd.n682 iovdd.n681 0.818682
R2939 iovdd.n680 iovdd.n623 0.818682
R2940 iovdd.n679 iovdd.n678 0.818682
R2941 iovdd.n625 iovdd.n624 0.818682
R2942 iovdd.n667 iovdd.n666 0.818682
R2943 iovdd.n665 iovdd.n632 0.818682
R2944 iovdd.n664 iovdd.n663 0.818682
R2945 iovdd.n634 iovdd.n633 0.818682
R2946 iovdd.n652 iovdd.n651 0.818682
R2947 iovdd.n650 iovdd.n641 0.818682
R2948 iovdd.n422 iovdd.n421 0.818682
R2949 iovdd.n1266 iovdd.n1265 0.818682
R2950 iovdd.n414 iovdd.n413 0.818682
R2951 iovdd.n1278 iovdd.n1277 0.818682
R2952 iovdd.n648 iovdd.n647 0.818682
R2953 iovdd.n643 iovdd.n641 0.818682
R2954 iovdd.n653 iovdd.n652 0.818682
R2955 iovdd.n654 iovdd.n634 0.818682
R2956 iovdd.n663 iovdd.n662 0.818682
R2957 iovdd.n636 iovdd.n632 0.818682
R2958 iovdd.n668 iovdd.n667 0.818682
R2959 iovdd.n669 iovdd.n625 0.818682
R2960 iovdd.n678 iovdd.n677 0.818682
R2961 iovdd.n627 iovdd.n623 0.818682
R2962 iovdd.n683 iovdd.n682 0.818682
R2963 iovdd.n684 iovdd.n616 0.818682
R2964 iovdd.n693 iovdd.n692 0.818682
R2965 iovdd.n618 iovdd.n614 0.818682
R2966 iovdd.n698 iovdd.n697 0.818682
R2967 iovdd.n699 iovdd.n607 0.818682
R2968 iovdd.n708 iovdd.n707 0.818682
R2969 iovdd.n609 iovdd.n605 0.818682
R2970 iovdd.n713 iovdd.n712 0.818682
R2971 iovdd.n714 iovdd.n598 0.818682
R2972 iovdd.n723 iovdd.n722 0.818682
R2973 iovdd.n600 iovdd.n596 0.818682
R2974 iovdd.n728 iovdd.n727 0.818682
R2975 iovdd.n729 iovdd.n589 0.818682
R2976 iovdd.n738 iovdd.n737 0.818682
R2977 iovdd.n591 iovdd.n587 0.818682
R2978 iovdd.n743 iovdd.n742 0.818682
R2979 iovdd.n744 iovdd.n580 0.818682
R2980 iovdd.n753 iovdd.n752 0.818682
R2981 iovdd.n582 iovdd.n578 0.818682
R2982 iovdd.n758 iovdd.n757 0.818682
R2983 iovdd.n759 iovdd.n571 0.818682
R2984 iovdd.n768 iovdd.n767 0.818682
R2985 iovdd.n573 iovdd.n421 0.818682
R2986 iovdd.n1267 iovdd.n1266 0.818682
R2987 iovdd.n1268 iovdd.n414 0.818682
R2988 iovdd.n1277 iovdd.n1276 0.818682
R2989 iovdd.n945 iovdd.n944 0.416993
R2990 iovdd.n650 iovdd.n649 0.416993
R2991 iovdd.n1239 iovdd 0.341436
R2992 iovdd.n939 iovdd.n937 0.201704
R2993 iovdd.n644 iovdd.n642 0.201704
R2994 iovdd.n1325 iovdd.n1324 0.2005
R2995 iovdd.n1317 iovdd.n242 0.2005
R2996 iovdd.n1320 iovdd.n1319 0.2005
R2997 iovdd.n245 iovdd.n244 0.2005
R2998 iovdd.n1061 iovdd.n1060 0.2005
R2999 iovdd.n869 iovdd.n867 0.2005
R3000 iovdd.n1056 iovdd.n1055 0.2005
R3001 iovdd.n872 iovdd.n871 0.2005
R3002 iovdd.n1046 iovdd.n1045 0.2005
R3003 iovdd.n878 iovdd.n876 0.2005
R3004 iovdd.n1041 iovdd.n1040 0.2005
R3005 iovdd.n881 iovdd.n880 0.2005
R3006 iovdd.n1031 iovdd.n1030 0.2005
R3007 iovdd.n887 iovdd.n885 0.2005
R3008 iovdd.n1026 iovdd.n1025 0.2005
R3009 iovdd.n890 iovdd.n889 0.2005
R3010 iovdd.n1016 iovdd.n1015 0.2005
R3011 iovdd.n896 iovdd.n894 0.2005
R3012 iovdd.n1011 iovdd.n1010 0.2005
R3013 iovdd.n899 iovdd.n898 0.2005
R3014 iovdd.n1001 iovdd.n1000 0.2005
R3015 iovdd.n905 iovdd.n903 0.2005
R3016 iovdd.n996 iovdd.n995 0.2005
R3017 iovdd.n908 iovdd.n907 0.2005
R3018 iovdd.n986 iovdd.n985 0.2005
R3019 iovdd.n914 iovdd.n912 0.2005
R3020 iovdd.n981 iovdd.n980 0.2005
R3021 iovdd.n917 iovdd.n916 0.2005
R3022 iovdd.n971 iovdd.n970 0.2005
R3023 iovdd.n923 iovdd.n921 0.2005
R3024 iovdd.n966 iovdd.n965 0.2005
R3025 iovdd.n926 iovdd.n925 0.2005
R3026 iovdd.n956 iovdd.n955 0.2005
R3027 iovdd.n932 iovdd.n930 0.2005
R3028 iovdd.n951 iovdd.n950 0.2005
R3029 iovdd.n935 iovdd.n934 0.2005
R3030 iovdd.n941 iovdd.n940 0.2005
R3031 iovdd.n1275 iovdd.n1274 0.2005
R3032 iovdd.n417 iovdd.n416 0.2005
R3033 iovdd.n1270 iovdd.n1269 0.2005
R3034 iovdd.n420 iovdd.n419 0.2005
R3035 iovdd.n766 iovdd.n765 0.2005
R3036 iovdd.n574 iovdd.n572 0.2005
R3037 iovdd.n761 iovdd.n760 0.2005
R3038 iovdd.n577 iovdd.n576 0.2005
R3039 iovdd.n751 iovdd.n750 0.2005
R3040 iovdd.n583 iovdd.n581 0.2005
R3041 iovdd.n746 iovdd.n745 0.2005
R3042 iovdd.n586 iovdd.n585 0.2005
R3043 iovdd.n736 iovdd.n735 0.2005
R3044 iovdd.n592 iovdd.n590 0.2005
R3045 iovdd.n731 iovdd.n730 0.2005
R3046 iovdd.n595 iovdd.n594 0.2005
R3047 iovdd.n721 iovdd.n720 0.2005
R3048 iovdd.n601 iovdd.n599 0.2005
R3049 iovdd.n716 iovdd.n715 0.2005
R3050 iovdd.n604 iovdd.n603 0.2005
R3051 iovdd.n706 iovdd.n705 0.2005
R3052 iovdd.n610 iovdd.n608 0.2005
R3053 iovdd.n701 iovdd.n700 0.2005
R3054 iovdd.n613 iovdd.n612 0.2005
R3055 iovdd.n691 iovdd.n690 0.2005
R3056 iovdd.n619 iovdd.n617 0.2005
R3057 iovdd.n686 iovdd.n685 0.2005
R3058 iovdd.n622 iovdd.n621 0.2005
R3059 iovdd.n676 iovdd.n675 0.2005
R3060 iovdd.n628 iovdd.n626 0.2005
R3061 iovdd.n671 iovdd.n670 0.2005
R3062 iovdd.n631 iovdd.n630 0.2005
R3063 iovdd.n661 iovdd.n660 0.2005
R3064 iovdd.n637 iovdd.n635 0.2005
R3065 iovdd.n656 iovdd.n655 0.2005
R3066 iovdd.n640 iovdd.n639 0.2005
R3067 iovdd.n646 iovdd.n645 0.2005
R3068 iovdd.n1357 iovdd 0.1105
R3069 iovdd.n275 iovdd 0.1105
R3070 iovdd.n1227 iovdd 0.1105
R3071 iovdd.n1324 iovdd.n1323 0.1105
R3072 iovdd.n1322 iovdd.n242 0.1105
R3073 iovdd.n1321 iovdd.n1320 0.1105
R3074 iovdd.n244 iovdd.n243 0.1105
R3075 iovdd.n1060 iovdd.n1059 0.1105
R3076 iovdd.n1058 iovdd.n869 0.1105
R3077 iovdd.n1057 iovdd.n1056 0.1105
R3078 iovdd.n871 iovdd.n870 0.1105
R3079 iovdd.n1045 iovdd.n1044 0.1105
R3080 iovdd.n1043 iovdd.n878 0.1105
R3081 iovdd.n1042 iovdd.n1041 0.1105
R3082 iovdd.n880 iovdd.n879 0.1105
R3083 iovdd.n1030 iovdd.n1029 0.1105
R3084 iovdd.n1028 iovdd.n887 0.1105
R3085 iovdd.n1027 iovdd.n1026 0.1105
R3086 iovdd.n889 iovdd.n888 0.1105
R3087 iovdd.n1015 iovdd.n1014 0.1105
R3088 iovdd.n1013 iovdd.n896 0.1105
R3089 iovdd.n1012 iovdd.n1011 0.1105
R3090 iovdd.n898 iovdd.n897 0.1105
R3091 iovdd.n1000 iovdd.n999 0.1105
R3092 iovdd.n998 iovdd.n905 0.1105
R3093 iovdd.n997 iovdd.n996 0.1105
R3094 iovdd.n907 iovdd.n906 0.1105
R3095 iovdd.n985 iovdd.n984 0.1105
R3096 iovdd.n983 iovdd.n914 0.1105
R3097 iovdd.n982 iovdd.n981 0.1105
R3098 iovdd.n916 iovdd.n915 0.1105
R3099 iovdd.n970 iovdd.n969 0.1105
R3100 iovdd.n968 iovdd.n923 0.1105
R3101 iovdd.n967 iovdd.n966 0.1105
R3102 iovdd.n925 iovdd.n924 0.1105
R3103 iovdd.n955 iovdd.n954 0.1105
R3104 iovdd.n953 iovdd.n932 0.1105
R3105 iovdd.n952 iovdd.n951 0.1105
R3106 iovdd.n934 iovdd.n933 0.1105
R3107 iovdd.n1274 iovdd.n1273 0.1105
R3108 iovdd.n1272 iovdd.n417 0.1105
R3109 iovdd.n1271 iovdd.n1270 0.1105
R3110 iovdd.n419 iovdd.n418 0.1105
R3111 iovdd.n765 iovdd.n764 0.1105
R3112 iovdd.n763 iovdd.n574 0.1105
R3113 iovdd.n762 iovdd.n761 0.1105
R3114 iovdd.n576 iovdd.n575 0.1105
R3115 iovdd.n750 iovdd.n749 0.1105
R3116 iovdd.n748 iovdd.n583 0.1105
R3117 iovdd.n747 iovdd.n746 0.1105
R3118 iovdd.n585 iovdd.n584 0.1105
R3119 iovdd.n735 iovdd.n734 0.1105
R3120 iovdd.n733 iovdd.n592 0.1105
R3121 iovdd.n732 iovdd.n731 0.1105
R3122 iovdd.n594 iovdd.n593 0.1105
R3123 iovdd.n720 iovdd.n719 0.1105
R3124 iovdd.n718 iovdd.n601 0.1105
R3125 iovdd.n717 iovdd.n716 0.1105
R3126 iovdd.n603 iovdd.n602 0.1105
R3127 iovdd.n705 iovdd.n704 0.1105
R3128 iovdd.n703 iovdd.n610 0.1105
R3129 iovdd.n702 iovdd.n701 0.1105
R3130 iovdd.n612 iovdd.n611 0.1105
R3131 iovdd.n690 iovdd.n689 0.1105
R3132 iovdd.n688 iovdd.n619 0.1105
R3133 iovdd.n687 iovdd.n686 0.1105
R3134 iovdd.n621 iovdd.n620 0.1105
R3135 iovdd.n675 iovdd.n674 0.1105
R3136 iovdd.n673 iovdd.n628 0.1105
R3137 iovdd.n672 iovdd.n671 0.1105
R3138 iovdd.n630 iovdd.n629 0.1105
R3139 iovdd.n660 iovdd.n659 0.1105
R3140 iovdd.n658 iovdd.n637 0.1105
R3141 iovdd.n657 iovdd.n656 0.1105
R3142 iovdd.n639 iovdd.n638 0.1105
R3143 iovdd.t0 iovdd.n8 0.063271
R3144 iovdd.t0 iovdd.n25 0.0625942
R3145 iovdd.t0 iovdd.n1360 0.0625838
R3146 iovdd.n1363 iovdd.n1 0.0607875
R3147 iovdd.n294 iovdd.n1 0.0607875
R3148 iovdd.n295 iovdd.n294 0.0607875
R3149 iovdd.n296 iovdd.n295 0.0607875
R3150 iovdd.n287 iovdd.n285 0.0607875
R3151 iovdd.n285 iovdd.n283 0.0607875
R3152 iovdd.n283 iovdd.n281 0.0607875
R3153 iovdd.n281 iovdd.n279 0.0607875
R3154 iovdd.n644 iovdd.n638 0.0568704
R3155 iovdd.n939 iovdd.n933 0.0568704
R3156 iovdd iovdd.n1363 0.041993
R3157 iovdd iovdd.n287 0.0350089
R3158 iovdd.n1294 iovdd.n1293 0.0347222
R3159 iovdd.n1293 iovdd.n1292 0.0347222
R3160 iovdd.n1292 iovdd.n1287 0.0347222
R3161 iovdd.n1287 iovdd.n1286 0.0347222
R3162 iovdd.n1188 iovdd.n1183 0.0347222
R3163 iovdd.n1189 iovdd.n1188 0.0347222
R3164 iovdd.n1190 iovdd.n1189 0.0347222
R3165 iovdd.n1190 iovdd.n1090 0.0347222
R3166 iovdd.n558 iovdd.n425 0.0347222
R3167 iovdd.n554 iovdd.n425 0.0347222
R3168 iovdd.n554 iovdd.n553 0.0347222
R3169 iovdd.n553 iovdd.n552 0.0347222
R3170 iovdd.n557 iovdd.n424 0.0347222
R3171 iovdd.n557 iovdd.n556 0.0347222
R3172 iovdd.n556 iovdd.n555 0.0347222
R3173 iovdd.n555 iovdd.n430 0.0347222
R3174 iovdd.n551 iovdd.n430 0.0347222
R3175 iovdd.n551 iovdd.n550 0.0347222
R3176 iovdd.n1185 iovdd.n771 0.0347222
R3177 iovdd.n1187 iovdd.n1185 0.0347222
R3178 iovdd.n1187 iovdd.n1182 0.0347222
R3179 iovdd.n1192 iovdd.n1182 0.0347222
R3180 iovdd.n1194 iovdd.n1192 0.0347222
R3181 iovdd.n1220 iovdd.n1194 0.0347222
R3182 iovdd.n1089 iovdd.n862 0.0347222
R3183 iovdd.n1226 iovdd.n862 0.0347222
R3184 iovdd.n1296 iovdd.n1295 0.0347222
R3185 iovdd.n1295 iovdd.n1285 0.0347222
R3186 iovdd.n1291 iovdd.n1285 0.0347222
R3187 iovdd.n1291 iovdd.n1290 0.0347222
R3188 iovdd.n1290 iovdd.n236 0.0347222
R3189 iovdd.n1354 iovdd.n236 0.0347222
R3190 iovdd.n212 iovdd.n80 0.0301825
R3191 iovdd.n524 iovdd.n330 0.0301825
R3192 iovdd.n1165 iovdd.n823 0.0301825
R3193 iovdd.n1228 iovdd.n858 0.0301825
R3194 iovdd.n45 iovdd.n44 0.0301825
R3195 iovdd.n403 iovdd.n54 0.0293095
R3196 iovdd.n125 iovdd.n71 0.0293095
R3197 iovdd.n143 iovdd.n88 0.0293095
R3198 iovdd.n159 iovdd.n105 0.0293095
R3199 iovdd.n1253 iovdd.n356 0.0293095
R3200 iovdd.n439 iovdd.n339 0.0293095
R3201 iovdd.n457 iovdd.n322 0.0293095
R3202 iovdd.n473 iovdd.n305 0.0293095
R3203 iovdd.n852 iovdd.n851 0.0293095
R3204 iovdd.n1097 iovdd.n831 0.0293095
R3205 iovdd.n1115 iovdd.n814 0.0293095
R3206 iovdd.n1131 iovdd.n797 0.0293095
R3207 iovdd.n133 iovdd.n79 0.0288977
R3208 iovdd.n447 iovdd.n331 0.0288977
R3209 iovdd.n1107 iovdd.n822 0.0288977
R3210 iovdd.n1289 iovdd.n62 0.0284365
R3211 iovdd.n238 iovdd.n63 0.0284365
R3212 iovdd.n188 iovdd.n96 0.0284365
R3213 iovdd.n185 iovdd.n97 0.0284365
R3214 iovdd.n429 iovdd.n348 0.0284365
R3215 iovdd.n549 iovdd.n347 0.0284365
R3216 iovdd.n500 iovdd.n314 0.0284365
R3217 iovdd.n497 iovdd.n313 0.0284365
R3218 iovdd.n1191 iovdd.n840 0.0284365
R3219 iovdd.n1219 iovdd.n839 0.0284365
R3220 iovdd.n1149 iovdd.n806 0.0284365
R3221 iovdd.n1147 iovdd.n805 0.0284365
R3222 iovdd.n1311 iovdd.n1310 0.0284365
R3223 iovdd.n290 iovdd.n277 0.0284365
R3224 iovdd.n399 iovdd.n55 0.0280247
R3225 iovdd.n227 iovdd.n70 0.0280247
R3226 iovdd.n197 iovdd.n89 0.0280247
R3227 iovdd.n176 iovdd.n104 0.0280247
R3228 iovdd.n1247 iovdd.n355 0.0280247
R3229 iovdd.n539 iovdd.n340 0.0280247
R3230 iovdd.n509 iovdd.n321 0.0280247
R3231 iovdd.n488 iovdd.n306 0.0280247
R3232 iovdd.n850 iovdd.n849 0.0280247
R3233 iovdd.n1175 iovdd.n832 0.0280247
R3234 iovdd.n1155 iovdd.n813 0.0280247
R3235 iovdd.n1141 iovdd.n798 0.0280247
R3236 iovdd.n406 iovdd.n53 0.0275635
R3237 iovdd.n127 iovdd.n72 0.0275635
R3238 iovdd.n141 iovdd.n87 0.0275635
R3239 iovdd.n161 iovdd.n106 0.0275635
R3240 iovdd.n1256 iovdd.n357 0.0275635
R3241 iovdd.n441 iovdd.n338 0.0275635
R3242 iovdd.n455 iovdd.n323 0.0275635
R3243 iovdd.n475 iovdd.n304 0.0275635
R3244 iovdd.n1231 iovdd.n1230 0.0275635
R3245 iovdd.n1099 iovdd.n830 0.0275635
R3246 iovdd.n1113 iovdd.n815 0.0275635
R3247 iovdd.n1133 iovdd.n796 0.0275635
R3248 iovdd.n1288 iovdd.n61 0.0271517
R3249 iovdd.n119 iovdd.n64 0.0271517
R3250 iovdd.n149 iovdd.n95 0.0271517
R3251 iovdd.n153 iovdd.n98 0.0271517
R3252 iovdd.n428 iovdd.n349 0.0271517
R3253 iovdd.n433 iovdd.n346 0.0271517
R3254 iovdd.n463 iovdd.n315 0.0271517
R3255 iovdd.n467 iovdd.n312 0.0271517
R3256 iovdd.n1181 iovdd.n841 0.0271517
R3257 iovdd.n1091 iovdd.n838 0.0271517
R3258 iovdd.n1121 iovdd.n807 0.0271517
R3259 iovdd.n1125 iovdd.n804 0.0271517
R3260 iovdd.n215 iovdd.n78 0.0266905
R3261 iovdd.n209 iovdd.n81 0.0266905
R3262 iovdd.n527 iovdd.n332 0.0266905
R3263 iovdd.n521 iovdd.n329 0.0266905
R3264 iovdd.n1167 iovdd.n824 0.0266905
R3265 iovdd.n1163 iovdd.n821 0.0266905
R3266 iovdd.n395 iovdd.n52 0.0262787
R3267 iovdd.n221 iovdd.n73 0.0262787
R3268 iovdd.n203 iovdd.n86 0.0262787
R3269 iovdd.n170 iovdd.n107 0.0262787
R3270 iovdd.n1243 iovdd.n358 0.0262787
R3271 iovdd.n533 iovdd.n337 0.0262787
R3272 iovdd.n515 iovdd.n324 0.0262787
R3273 iovdd.n482 iovdd.n303 0.0262787
R3274 iovdd.n853 iovdd.n790 0.0262787
R3275 iovdd.n1171 iovdd.n829 0.0262787
R3276 iovdd.n1159 iovdd.n816 0.0262787
R3277 iovdd.n1137 iovdd.n795 0.0262787
R3278 iovdd.n1299 iovdd.n56 0.0258175
R3279 iovdd.n123 iovdd.n69 0.0258175
R3280 iovdd.n145 iovdd.n90 0.0258175
R3281 iovdd.n157 iovdd.n103 0.0258175
R3282 iovdd.n1250 iovdd.n354 0.0258175
R3283 iovdd.n437 iovdd.n341 0.0258175
R3284 iovdd.n459 iovdd.n320 0.0258175
R3285 iovdd.n471 iovdd.n307 0.0258175
R3286 iovdd.n848 iovdd.n847 0.0258175
R3287 iovdd.n1095 iovdd.n833 0.0258175
R3288 iovdd.n1117 iovdd.n812 0.0258175
R3289 iovdd.n1129 iovdd.n799 0.0258175
R3290 iovdd.n131 iovdd.n77 0.0254057
R3291 iovdd.n137 iovdd.n82 0.0254057
R3292 iovdd.n445 iovdd.n333 0.0254057
R3293 iovdd.n451 iovdd.n328 0.0254057
R3294 iovdd.n1103 iovdd.n825 0.0254057
R3295 iovdd.n1109 iovdd.n820 0.0254057
R3296 iovdd.n1284 iovdd.n60 0.0249444
R3297 iovdd.n233 iovdd.n65 0.0249444
R3298 iovdd.n191 iovdd.n94 0.0249444
R3299 iovdd.n182 iovdd.n99 0.0249444
R3300 iovdd.n427 iovdd.n350 0.0249444
R3301 iovdd.n545 iovdd.n345 0.0249444
R3302 iovdd.n503 iovdd.n316 0.0249444
R3303 iovdd.n494 iovdd.n311 0.0249444
R3304 iovdd.n1186 iovdd.n842 0.0249444
R3305 iovdd.n1179 iovdd.n837 0.0249444
R3306 iovdd.n1151 iovdd.n808 0.0249444
R3307 iovdd.n1145 iovdd.n803 0.0249444
R3308 iovdd.n1282 iovdd.n57 0.0245327
R3309 iovdd.n230 iovdd.n68 0.0245327
R3310 iovdd.n194 iovdd.n91 0.0245327
R3311 iovdd.n179 iovdd.n102 0.0245327
R3312 iovdd.n423 iovdd.n353 0.0245327
R3313 iovdd.n542 iovdd.n342 0.0245327
R3314 iovdd.n506 iovdd.n319 0.0245327
R3315 iovdd.n491 iovdd.n308 0.0245327
R3316 iovdd.n846 iovdd.n845 0.0245327
R3317 iovdd.n1177 iovdd.n834 0.0245327
R3318 iovdd.n1153 iovdd.n811 0.0245327
R3319 iovdd.n1143 iovdd.n800 0.0245327
R3320 iovdd.n279 iovdd.n111 0.0245327
R3321 iovdd.n409 iovdd.n51 0.0240714
R3322 iovdd.n129 iovdd.n74 0.0240714
R3323 iovdd.n139 iovdd.n85 0.0240714
R3324 iovdd.n163 iovdd.n108 0.0240714
R3325 iovdd.n1259 iovdd.n359 0.0240714
R3326 iovdd.n443 iovdd.n336 0.0240714
R3327 iovdd.n453 iovdd.n325 0.0240714
R3328 iovdd.n478 iovdd.n302 0.0240714
R3329 iovdd.n854 iovdd.n780 0.0240714
R3330 iovdd.n1101 iovdd.n828 0.0240714
R3331 iovdd.n1111 iovdd.n817 0.0240714
R3332 iovdd.n1135 iovdd.n794 0.0240714
R3333 iovdd.n1283 iovdd.n59 0.0236596
R3334 iovdd.n121 iovdd.n66 0.0236596
R3335 iovdd.n147 iovdd.n93 0.0236596
R3336 iovdd.n155 iovdd.n100 0.0236596
R3337 iovdd.n426 iovdd.n351 0.0236596
R3338 iovdd.n435 iovdd.n344 0.0236596
R3339 iovdd.n461 iovdd.n317 0.0236596
R3340 iovdd.n469 iovdd.n310 0.0236596
R3341 iovdd.n1184 iovdd.n843 0.0236596
R3342 iovdd.n1093 iovdd.n836 0.0236596
R3343 iovdd.n1119 iovdd.n809 0.0236596
R3344 iovdd.n1127 iovdd.n802 0.0236596
R3345 iovdd.n393 iovdd.n46 0.0231984
R3346 iovdd.n218 iovdd.n76 0.0231984
R3347 iovdd.n206 iovdd.n83 0.0231984
R3348 iovdd.n167 iovdd.n110 0.0231984
R3349 iovdd.n1241 iovdd.n361 0.0231984
R3350 iovdd.n530 iovdd.n334 0.0231984
R3351 iovdd.n518 iovdd.n327 0.0231984
R3352 iovdd.n300 iovdd.n299 0.0231984
R3353 iovdd.n855 iovdd.n567 0.0231984
R3354 iovdd.n1169 iovdd.n826 0.0231984
R3355 iovdd.n1161 iovdd.n819 0.0231984
R3356 iovdd.n1088 iovdd.n792 0.0231984
R3357 iovdd.n393 iovdd.n50 0.0227866
R3358 iovdd.n218 iovdd.n75 0.0227866
R3359 iovdd.n206 iovdd.n84 0.0227866
R3360 iovdd.n167 iovdd.n109 0.0227866
R3361 iovdd.n1241 iovdd.n360 0.0227866
R3362 iovdd.n530 iovdd.n335 0.0227866
R3363 iovdd.n518 iovdd.n326 0.0227866
R3364 iovdd.n301 iovdd.n300 0.0227866
R3365 iovdd.n856 iovdd.n855 0.0227866
R3366 iovdd.n1169 iovdd.n827 0.0227866
R3367 iovdd.n1161 iovdd.n818 0.0227866
R3368 iovdd.n1088 iovdd.n793 0.0227866
R3369 iovdd.n1283 iovdd.n58 0.0223254
R3370 iovdd.n121 iovdd.n67 0.0223254
R3371 iovdd.n147 iovdd.n92 0.0223254
R3372 iovdd.n155 iovdd.n101 0.0223254
R3373 iovdd.n426 iovdd.n352 0.0223254
R3374 iovdd.n435 iovdd.n343 0.0223254
R3375 iovdd.n461 iovdd.n318 0.0223254
R3376 iovdd.n469 iovdd.n309 0.0223254
R3377 iovdd.n1184 iovdd.n844 0.0223254
R3378 iovdd.n1093 iovdd.n835 0.0223254
R3379 iovdd.n1119 iovdd.n810 0.0223254
R3380 iovdd.n1127 iovdd.n801 0.0223254
R3381 iovdd.n1227 iovdd.n861 0.0223254
R3382 iovdd.n1358 iovdd.n1357 0.0223254
R3383 iovdd.n409 iovdd.n50 0.0219136
R3384 iovdd.n129 iovdd.n75 0.0219136
R3385 iovdd.n139 iovdd.n84 0.0219136
R3386 iovdd.n163 iovdd.n109 0.0219136
R3387 iovdd.n1259 iovdd.n360 0.0219136
R3388 iovdd.n443 iovdd.n335 0.0219136
R3389 iovdd.n453 iovdd.n326 0.0219136
R3390 iovdd.n478 iovdd.n301 0.0219136
R3391 iovdd.n856 iovdd.n780 0.0219136
R3392 iovdd.n1101 iovdd.n827 0.0219136
R3393 iovdd.n1111 iovdd.n818 0.0219136
R3394 iovdd.n1135 iovdd.n793 0.0219136
R3395 iovdd.n1282 iovdd.n58 0.0214524
R3396 iovdd.n230 iovdd.n67 0.0214524
R3397 iovdd.n194 iovdd.n92 0.0214524
R3398 iovdd.n179 iovdd.n101 0.0214524
R3399 iovdd.n423 iovdd.n352 0.0214524
R3400 iovdd.n542 iovdd.n343 0.0214524
R3401 iovdd.n506 iovdd.n318 0.0214524
R3402 iovdd.n491 iovdd.n309 0.0214524
R3403 iovdd.n845 iovdd.n844 0.0214524
R3404 iovdd.n1177 iovdd.n835 0.0214524
R3405 iovdd.n1153 iovdd.n810 0.0214524
R3406 iovdd.n1143 iovdd.n801 0.0214524
R3407 iovdd.n1225 iovdd.n861 0.0214524
R3408 iovdd.n1358 iovdd.n111 0.0214524
R3409 iovdd.n1284 iovdd.n59 0.0210406
R3410 iovdd.n233 iovdd.n66 0.0210406
R3411 iovdd.n191 iovdd.n93 0.0210406
R3412 iovdd.n182 iovdd.n100 0.0210406
R3413 iovdd.n427 iovdd.n351 0.0210406
R3414 iovdd.n545 iovdd.n344 0.0210406
R3415 iovdd.n503 iovdd.n317 0.0210406
R3416 iovdd.n494 iovdd.n310 0.0210406
R3417 iovdd.n1186 iovdd.n843 0.0210406
R3418 iovdd.n1179 iovdd.n836 0.0210406
R3419 iovdd.n1151 iovdd.n809 0.0210406
R3420 iovdd.n1145 iovdd.n802 0.0210406
R3421 iovdd.n412 iovdd.n46 0.0205794
R3422 iovdd.n131 iovdd.n76 0.0205794
R3423 iovdd.n137 iovdd.n83 0.0205794
R3424 iovdd.n112 iovdd.n110 0.0205794
R3425 iovdd.n1240 iovdd.n361 0.0205794
R3426 iovdd.n445 iovdd.n334 0.0205794
R3427 iovdd.n451 iovdd.n327 0.0205794
R3428 iovdd.n299 iovdd.n298 0.0205794
R3429 iovdd.n1238 iovdd.n567 0.0205794
R3430 iovdd.n1103 iovdd.n826 0.0205794
R3431 iovdd.n1109 iovdd.n819 0.0205794
R3432 iovdd.n859 iovdd.n792 0.0205794
R3433 iovdd.n1299 iovdd.n57 0.0201676
R3434 iovdd.n123 iovdd.n68 0.0201676
R3435 iovdd.n145 iovdd.n91 0.0201676
R3436 iovdd.n157 iovdd.n102 0.0201676
R3437 iovdd.n1250 iovdd.n353 0.0201676
R3438 iovdd.n437 iovdd.n342 0.0201676
R3439 iovdd.n459 iovdd.n319 0.0201676
R3440 iovdd.n471 iovdd.n308 0.0201676
R3441 iovdd.n847 iovdd.n846 0.0201676
R3442 iovdd.n1095 iovdd.n834 0.0201676
R3443 iovdd.n1117 iovdd.n811 0.0201676
R3444 iovdd.n1129 iovdd.n800 0.0201676
R3445 iovdd.n395 iovdd.n51 0.0197063
R3446 iovdd.n221 iovdd.n74 0.0197063
R3447 iovdd.n203 iovdd.n85 0.0197063
R3448 iovdd.n170 iovdd.n108 0.0197063
R3449 iovdd.n1243 iovdd.n359 0.0197063
R3450 iovdd.n533 iovdd.n336 0.0197063
R3451 iovdd.n515 iovdd.n325 0.0197063
R3452 iovdd.n482 iovdd.n302 0.0197063
R3453 iovdd.n854 iovdd.n853 0.0197063
R3454 iovdd.n1171 iovdd.n828 0.0197063
R3455 iovdd.n1159 iovdd.n817 0.0197063
R3456 iovdd.n1137 iovdd.n794 0.0197063
R3457 iovdd.n215 iovdd.n77 0.0192946
R3458 iovdd.n209 iovdd.n82 0.0192946
R3459 iovdd.n527 iovdd.n333 0.0192946
R3460 iovdd.n521 iovdd.n328 0.0192946
R3461 iovdd.n1167 iovdd.n825 0.0192946
R3462 iovdd.n1163 iovdd.n820 0.0192946
R3463 iovdd.n1288 iovdd.n60 0.0188333
R3464 iovdd.n119 iovdd.n65 0.0188333
R3465 iovdd.n149 iovdd.n94 0.0188333
R3466 iovdd.n153 iovdd.n99 0.0188333
R3467 iovdd.n428 iovdd.n350 0.0188333
R3468 iovdd.n433 iovdd.n345 0.0188333
R3469 iovdd.n463 iovdd.n316 0.0188333
R3470 iovdd.n467 iovdd.n311 0.0188333
R3471 iovdd.n1181 iovdd.n842 0.0188333
R3472 iovdd.n1091 iovdd.n837 0.0188333
R3473 iovdd.n1121 iovdd.n808 0.0188333
R3474 iovdd.n1125 iovdd.n803 0.0188333
R3475 iovdd.n406 iovdd.n52 0.0184215
R3476 iovdd.n127 iovdd.n73 0.0184215
R3477 iovdd.n141 iovdd.n86 0.0184215
R3478 iovdd.n161 iovdd.n107 0.0184215
R3479 iovdd.n1256 iovdd.n358 0.0184215
R3480 iovdd.n441 iovdd.n337 0.0184215
R3481 iovdd.n455 iovdd.n324 0.0184215
R3482 iovdd.n475 iovdd.n303 0.0184215
R3483 iovdd.n1231 iovdd.n790 0.0184215
R3484 iovdd.n1099 iovdd.n829 0.0184215
R3485 iovdd.n1113 iovdd.n816 0.0184215
R3486 iovdd.n1133 iovdd.n795 0.0184215
R3487 iovdd.n565 iovdd.n564 0.0180786
R3488 iovdd.n1263 iovdd.n1262 0.0180786
R3489 iovdd.n1242 iovdd.n566 0.0180786
R3490 iovdd.n1260 iovdd.n563 0.0180786
R3491 iovdd.n1258 iovdd.n1244 0.0180786
R3492 iovdd.n1257 iovdd.n562 0.0180786
R3493 iovdd.n1255 iovdd.n1246 0.0180786
R3494 iovdd.n1254 iovdd.n561 0.0180786
R3495 iovdd.n1252 iovdd.n1248 0.0180786
R3496 iovdd.n1251 iovdd.n560 0.0180786
R3497 iovdd.n1249 iovdd.n424 0.0180786
R3498 iovdd.n434 iovdd.n249 0.0180786
R3499 iovdd.n546 iovdd.n544 0.0180786
R3500 iovdd.n436 iovdd.n250 0.0180786
R3501 iovdd.n543 iovdd.n541 0.0180786
R3502 iovdd.n438 iovdd.n251 0.0180786
R3503 iovdd.n540 iovdd.n538 0.0180786
R3504 iovdd.n440 iovdd.n252 0.0180786
R3505 iovdd.n537 iovdd.n535 0.0180786
R3506 iovdd.n442 iovdd.n253 0.0180786
R3507 iovdd.n534 iovdd.n532 0.0180786
R3508 iovdd.n444 iovdd.n254 0.0180786
R3509 iovdd.n531 iovdd.n529 0.0180786
R3510 iovdd.n446 iovdd.n255 0.0180786
R3511 iovdd.n528 iovdd.n526 0.0180786
R3512 iovdd.n448 iovdd.n256 0.0180786
R3513 iovdd.n525 iovdd.n523 0.0180786
R3514 iovdd.n450 iovdd.n257 0.0180786
R3515 iovdd.n522 iovdd.n520 0.0180786
R3516 iovdd.n452 iovdd.n258 0.0180786
R3517 iovdd.n519 iovdd.n517 0.0180786
R3518 iovdd.n454 iovdd.n259 0.0180786
R3519 iovdd.n516 iovdd.n514 0.0180786
R3520 iovdd.n456 iovdd.n260 0.0180786
R3521 iovdd.n513 iovdd.n511 0.0180786
R3522 iovdd.n458 iovdd.n261 0.0180786
R3523 iovdd.n510 iovdd.n508 0.0180786
R3524 iovdd.n460 iovdd.n262 0.0180786
R3525 iovdd.n507 iovdd.n505 0.0180786
R3526 iovdd.n462 iovdd.n263 0.0180786
R3527 iovdd.n504 iovdd.n502 0.0180786
R3528 iovdd.n464 iovdd.n264 0.0180786
R3529 iovdd.n501 iovdd.n499 0.0180786
R3530 iovdd.n466 iovdd.n265 0.0180786
R3531 iovdd.n498 iovdd.n496 0.0180786
R3532 iovdd.n468 iovdd.n266 0.0180786
R3533 iovdd.n495 iovdd.n493 0.0180786
R3534 iovdd.n470 iovdd.n267 0.0180786
R3535 iovdd.n492 iovdd.n490 0.0180786
R3536 iovdd.n472 iovdd.n268 0.0180786
R3537 iovdd.n489 iovdd.n487 0.0180786
R3538 iovdd.n474 iovdd.n269 0.0180786
R3539 iovdd.n486 iovdd.n484 0.0180786
R3540 iovdd.n476 iovdd.n270 0.0180786
R3541 iovdd.n483 iovdd.n481 0.0180786
R3542 iovdd.n479 iovdd.n271 0.0180786
R3543 iovdd.n477 iovdd.n273 0.0180786
R3544 iovdd.n480 iovdd.n272 0.0180786
R3545 iovdd.n1312 iovdd.n274 0.0180786
R3546 iovdd.n1312 iovdd.n276 0.0180786
R3547 iovdd.n274 iovdd.n272 0.0180786
R3548 iovdd.n480 iovdd.n273 0.0180786
R3549 iovdd.n479 iovdd.n477 0.0180786
R3550 iovdd.n483 iovdd.n271 0.0180786
R3551 iovdd.n481 iovdd.n476 0.0180786
R3552 iovdd.n486 iovdd.n270 0.0180786
R3553 iovdd.n484 iovdd.n474 0.0180786
R3554 iovdd.n489 iovdd.n269 0.0180786
R3555 iovdd.n487 iovdd.n472 0.0180786
R3556 iovdd.n492 iovdd.n268 0.0180786
R3557 iovdd.n490 iovdd.n470 0.0180786
R3558 iovdd.n495 iovdd.n267 0.0180786
R3559 iovdd.n493 iovdd.n468 0.0180786
R3560 iovdd.n498 iovdd.n266 0.0180786
R3561 iovdd.n496 iovdd.n466 0.0180786
R3562 iovdd.n501 iovdd.n265 0.0180786
R3563 iovdd.n499 iovdd.n464 0.0180786
R3564 iovdd.n504 iovdd.n264 0.0180786
R3565 iovdd.n502 iovdd.n462 0.0180786
R3566 iovdd.n507 iovdd.n263 0.0180786
R3567 iovdd.n505 iovdd.n460 0.0180786
R3568 iovdd.n510 iovdd.n262 0.0180786
R3569 iovdd.n508 iovdd.n458 0.0180786
R3570 iovdd.n513 iovdd.n261 0.0180786
R3571 iovdd.n511 iovdd.n456 0.0180786
R3572 iovdd.n516 iovdd.n260 0.0180786
R3573 iovdd.n514 iovdd.n454 0.0180786
R3574 iovdd.n519 iovdd.n259 0.0180786
R3575 iovdd.n517 iovdd.n452 0.0180786
R3576 iovdd.n522 iovdd.n258 0.0180786
R3577 iovdd.n520 iovdd.n450 0.0180786
R3578 iovdd.n525 iovdd.n257 0.0180786
R3579 iovdd.n523 iovdd.n448 0.0180786
R3580 iovdd.n528 iovdd.n256 0.0180786
R3581 iovdd.n526 iovdd.n446 0.0180786
R3582 iovdd.n531 iovdd.n255 0.0180786
R3583 iovdd.n529 iovdd.n444 0.0180786
R3584 iovdd.n534 iovdd.n254 0.0180786
R3585 iovdd.n532 iovdd.n442 0.0180786
R3586 iovdd.n537 iovdd.n253 0.0180786
R3587 iovdd.n535 iovdd.n440 0.0180786
R3588 iovdd.n540 iovdd.n252 0.0180786
R3589 iovdd.n538 iovdd.n438 0.0180786
R3590 iovdd.n543 iovdd.n251 0.0180786
R3591 iovdd.n541 iovdd.n436 0.0180786
R3592 iovdd.n546 iovdd.n250 0.0180786
R3593 iovdd.n544 iovdd.n434 0.0180786
R3594 iovdd.n550 iovdd.n249 0.0180786
R3595 iovdd.n297 iovdd.n276 0.0180786
R3596 iovdd.n773 iovdd.n770 0.0180786
R3597 iovdd.n1237 iovdd.n568 0.0180786
R3598 iovdd.n778 iovdd.n569 0.0180786
R3599 iovdd.n1235 iovdd.n1234 0.0180786
R3600 iovdd.n782 iovdd.n779 0.0180786
R3601 iovdd.n1232 iovdd.n777 0.0180786
R3602 iovdd.n789 iovdd.n783 0.0180786
R3603 iovdd.n788 iovdd.n776 0.0180786
R3604 iovdd.n787 iovdd.n784 0.0180786
R3605 iovdd.n786 iovdd.n775 0.0180786
R3606 iovdd.n785 iovdd.n771 0.0180786
R3607 iovdd.n1220 iovdd.n1065 0.0180786
R3608 iovdd.n1195 iovdd.n1092 0.0180786
R3609 iovdd.n1180 iovdd.n1066 0.0180786
R3610 iovdd.n1196 iovdd.n1094 0.0180786
R3611 iovdd.n1178 iovdd.n1067 0.0180786
R3612 iovdd.n1197 iovdd.n1096 0.0180786
R3613 iovdd.n1176 iovdd.n1068 0.0180786
R3614 iovdd.n1198 iovdd.n1098 0.0180786
R3615 iovdd.n1174 iovdd.n1069 0.0180786
R3616 iovdd.n1199 iovdd.n1100 0.0180786
R3617 iovdd.n1172 iovdd.n1070 0.0180786
R3618 iovdd.n1200 iovdd.n1102 0.0180786
R3619 iovdd.n1170 iovdd.n1071 0.0180786
R3620 iovdd.n1201 iovdd.n1104 0.0180786
R3621 iovdd.n1168 iovdd.n1072 0.0180786
R3622 iovdd.n1202 iovdd.n1106 0.0180786
R3623 iovdd.n1166 iovdd.n1073 0.0180786
R3624 iovdd.n1203 iovdd.n1108 0.0180786
R3625 iovdd.n1164 iovdd.n1074 0.0180786
R3626 iovdd.n1204 iovdd.n1110 0.0180786
R3627 iovdd.n1162 iovdd.n1075 0.0180786
R3628 iovdd.n1205 iovdd.n1112 0.0180786
R3629 iovdd.n1160 iovdd.n1076 0.0180786
R3630 iovdd.n1206 iovdd.n1114 0.0180786
R3631 iovdd.n1158 iovdd.n1077 0.0180786
R3632 iovdd.n1207 iovdd.n1116 0.0180786
R3633 iovdd.n1156 iovdd.n1078 0.0180786
R3634 iovdd.n1208 iovdd.n1118 0.0180786
R3635 iovdd.n1154 iovdd.n1079 0.0180786
R3636 iovdd.n1209 iovdd.n1120 0.0180786
R3637 iovdd.n1152 iovdd.n1080 0.0180786
R3638 iovdd.n1210 iovdd.n1122 0.0180786
R3639 iovdd.n1150 iovdd.n1081 0.0180786
R3640 iovdd.n1211 iovdd.n1124 0.0180786
R3641 iovdd.n1148 iovdd.n1082 0.0180786
R3642 iovdd.n1212 iovdd.n1126 0.0180786
R3643 iovdd.n1146 iovdd.n1083 0.0180786
R3644 iovdd.n1213 iovdd.n1128 0.0180786
R3645 iovdd.n1144 iovdd.n1084 0.0180786
R3646 iovdd.n1214 iovdd.n1130 0.0180786
R3647 iovdd.n1142 iovdd.n1085 0.0180786
R3648 iovdd.n1215 iovdd.n1132 0.0180786
R3649 iovdd.n1140 iovdd.n1086 0.0180786
R3650 iovdd.n1216 iovdd.n1134 0.0180786
R3651 iovdd.n1138 iovdd.n1087 0.0180786
R3652 iovdd.n1217 iovdd.n1136 0.0180786
R3653 iovdd.n1226 iovdd.n1224 0.0180786
R3654 iovdd.n1217 iovdd.n1089 0.0180786
R3655 iovdd.n1136 iovdd.n1087 0.0180786
R3656 iovdd.n1216 iovdd.n1138 0.0180786
R3657 iovdd.n1134 iovdd.n1086 0.0180786
R3658 iovdd.n1215 iovdd.n1140 0.0180786
R3659 iovdd.n1132 iovdd.n1085 0.0180786
R3660 iovdd.n1214 iovdd.n1142 0.0180786
R3661 iovdd.n1130 iovdd.n1084 0.0180786
R3662 iovdd.n1213 iovdd.n1144 0.0180786
R3663 iovdd.n1128 iovdd.n1083 0.0180786
R3664 iovdd.n1212 iovdd.n1146 0.0180786
R3665 iovdd.n1126 iovdd.n1082 0.0180786
R3666 iovdd.n1211 iovdd.n1148 0.0180786
R3667 iovdd.n1124 iovdd.n1081 0.0180786
R3668 iovdd.n1210 iovdd.n1150 0.0180786
R3669 iovdd.n1122 iovdd.n1080 0.0180786
R3670 iovdd.n1209 iovdd.n1152 0.0180786
R3671 iovdd.n1120 iovdd.n1079 0.0180786
R3672 iovdd.n1208 iovdd.n1154 0.0180786
R3673 iovdd.n1118 iovdd.n1078 0.0180786
R3674 iovdd.n1207 iovdd.n1156 0.0180786
R3675 iovdd.n1116 iovdd.n1077 0.0180786
R3676 iovdd.n1206 iovdd.n1158 0.0180786
R3677 iovdd.n1114 iovdd.n1076 0.0180786
R3678 iovdd.n1205 iovdd.n1160 0.0180786
R3679 iovdd.n1112 iovdd.n1075 0.0180786
R3680 iovdd.n1204 iovdd.n1162 0.0180786
R3681 iovdd.n1110 iovdd.n1074 0.0180786
R3682 iovdd.n1203 iovdd.n1164 0.0180786
R3683 iovdd.n1108 iovdd.n1073 0.0180786
R3684 iovdd.n1202 iovdd.n1166 0.0180786
R3685 iovdd.n1106 iovdd.n1072 0.0180786
R3686 iovdd.n1201 iovdd.n1168 0.0180786
R3687 iovdd.n1104 iovdd.n1071 0.0180786
R3688 iovdd.n1200 iovdd.n1170 0.0180786
R3689 iovdd.n1102 iovdd.n1070 0.0180786
R3690 iovdd.n1199 iovdd.n1172 0.0180786
R3691 iovdd.n1100 iovdd.n1069 0.0180786
R3692 iovdd.n1198 iovdd.n1174 0.0180786
R3693 iovdd.n1098 iovdd.n1068 0.0180786
R3694 iovdd.n1197 iovdd.n1176 0.0180786
R3695 iovdd.n1096 iovdd.n1067 0.0180786
R3696 iovdd.n1196 iovdd.n1178 0.0180786
R3697 iovdd.n1094 iovdd.n1066 0.0180786
R3698 iovdd.n1195 iovdd.n1180 0.0180786
R3699 iovdd.n1092 iovdd.n1065 0.0180786
R3700 iovdd.n1224 iovdd.n860 0.0180786
R3701 iovdd.n392 iovdd.n390 0.0180786
R3702 iovdd.n1303 iovdd.n411 0.0180786
R3703 iovdd.n1302 iovdd.n394 0.0180786
R3704 iovdd.n410 iovdd.n408 0.0180786
R3705 iovdd.n1279 iovdd.n396 0.0180786
R3706 iovdd.n407 iovdd.n405 0.0180786
R3707 iovdd.n1280 iovdd.n398 0.0180786
R3708 iovdd.n404 iovdd.n402 0.0180786
R3709 iovdd.n1281 iovdd.n400 0.0180786
R3710 iovdd.n1300 iovdd.n1298 0.0180786
R3711 iovdd.n1296 iovdd.n401 0.0180786
R3712 iovdd.n237 iovdd.n120 0.0180786
R3713 iovdd.n1352 iovdd.n234 0.0180786
R3714 iovdd.n232 iovdd.n122 0.0180786
R3715 iovdd.n1351 iovdd.n231 0.0180786
R3716 iovdd.n229 iovdd.n124 0.0180786
R3717 iovdd.n1350 iovdd.n228 0.0180786
R3718 iovdd.n226 iovdd.n126 0.0180786
R3719 iovdd.n1349 iovdd.n225 0.0180786
R3720 iovdd.n223 iovdd.n128 0.0180786
R3721 iovdd.n1348 iovdd.n222 0.0180786
R3722 iovdd.n220 iovdd.n130 0.0180786
R3723 iovdd.n1347 iovdd.n219 0.0180786
R3724 iovdd.n217 iovdd.n132 0.0180786
R3725 iovdd.n1346 iovdd.n216 0.0180786
R3726 iovdd.n214 iovdd.n134 0.0180786
R3727 iovdd.n1345 iovdd.n213 0.0180786
R3728 iovdd.n211 iovdd.n136 0.0180786
R3729 iovdd.n1344 iovdd.n210 0.0180786
R3730 iovdd.n208 iovdd.n138 0.0180786
R3731 iovdd.n1343 iovdd.n207 0.0180786
R3732 iovdd.n205 iovdd.n140 0.0180786
R3733 iovdd.n1342 iovdd.n204 0.0180786
R3734 iovdd.n202 iovdd.n142 0.0180786
R3735 iovdd.n1341 iovdd.n201 0.0180786
R3736 iovdd.n199 iovdd.n144 0.0180786
R3737 iovdd.n1340 iovdd.n198 0.0180786
R3738 iovdd.n196 iovdd.n146 0.0180786
R3739 iovdd.n1339 iovdd.n195 0.0180786
R3740 iovdd.n193 iovdd.n148 0.0180786
R3741 iovdd.n1338 iovdd.n192 0.0180786
R3742 iovdd.n190 iovdd.n150 0.0180786
R3743 iovdd.n1337 iovdd.n189 0.0180786
R3744 iovdd.n187 iovdd.n152 0.0180786
R3745 iovdd.n1336 iovdd.n186 0.0180786
R3746 iovdd.n184 iovdd.n154 0.0180786
R3747 iovdd.n1335 iovdd.n183 0.0180786
R3748 iovdd.n181 iovdd.n156 0.0180786
R3749 iovdd.n1334 iovdd.n180 0.0180786
R3750 iovdd.n178 iovdd.n158 0.0180786
R3751 iovdd.n1333 iovdd.n177 0.0180786
R3752 iovdd.n175 iovdd.n160 0.0180786
R3753 iovdd.n1332 iovdd.n174 0.0180786
R3754 iovdd.n172 iovdd.n162 0.0180786
R3755 iovdd.n1331 iovdd.n171 0.0180786
R3756 iovdd.n169 iovdd.n164 0.0180786
R3757 iovdd.n1330 iovdd.n168 0.0180786
R3758 iovdd.n166 iovdd.n165 0.0180786
R3759 iovdd.n165 iovdd.n114 0.0180786
R3760 iovdd.n1356 iovdd.n117 0.0180786
R3761 iovdd.n117 iovdd.n113 0.0180786
R3762 iovdd.n168 iovdd.n166 0.0180786
R3763 iovdd.n1330 iovdd.n164 0.0180786
R3764 iovdd.n171 iovdd.n169 0.0180786
R3765 iovdd.n1331 iovdd.n162 0.0180786
R3766 iovdd.n174 iovdd.n172 0.0180786
R3767 iovdd.n1332 iovdd.n160 0.0180786
R3768 iovdd.n177 iovdd.n175 0.0180786
R3769 iovdd.n1333 iovdd.n158 0.0180786
R3770 iovdd.n180 iovdd.n178 0.0180786
R3771 iovdd.n1334 iovdd.n156 0.0180786
R3772 iovdd.n183 iovdd.n181 0.0180786
R3773 iovdd.n1335 iovdd.n154 0.0180786
R3774 iovdd.n186 iovdd.n184 0.0180786
R3775 iovdd.n1336 iovdd.n152 0.0180786
R3776 iovdd.n189 iovdd.n187 0.0180786
R3777 iovdd.n1337 iovdd.n150 0.0180786
R3778 iovdd.n192 iovdd.n190 0.0180786
R3779 iovdd.n1338 iovdd.n148 0.0180786
R3780 iovdd.n195 iovdd.n193 0.0180786
R3781 iovdd.n1339 iovdd.n146 0.0180786
R3782 iovdd.n198 iovdd.n196 0.0180786
R3783 iovdd.n1340 iovdd.n144 0.0180786
R3784 iovdd.n201 iovdd.n199 0.0180786
R3785 iovdd.n1341 iovdd.n142 0.0180786
R3786 iovdd.n204 iovdd.n202 0.0180786
R3787 iovdd.n1342 iovdd.n140 0.0180786
R3788 iovdd.n207 iovdd.n205 0.0180786
R3789 iovdd.n1343 iovdd.n138 0.0180786
R3790 iovdd.n210 iovdd.n208 0.0180786
R3791 iovdd.n1344 iovdd.n136 0.0180786
R3792 iovdd.n213 iovdd.n211 0.0180786
R3793 iovdd.n1345 iovdd.n134 0.0180786
R3794 iovdd.n216 iovdd.n214 0.0180786
R3795 iovdd.n1346 iovdd.n132 0.0180786
R3796 iovdd.n219 iovdd.n217 0.0180786
R3797 iovdd.n1347 iovdd.n130 0.0180786
R3798 iovdd.n222 iovdd.n220 0.0180786
R3799 iovdd.n1348 iovdd.n128 0.0180786
R3800 iovdd.n225 iovdd.n223 0.0180786
R3801 iovdd.n1349 iovdd.n126 0.0180786
R3802 iovdd.n228 iovdd.n226 0.0180786
R3803 iovdd.n1350 iovdd.n124 0.0180786
R3804 iovdd.n231 iovdd.n229 0.0180786
R3805 iovdd.n1351 iovdd.n122 0.0180786
R3806 iovdd.n234 iovdd.n232 0.0180786
R3807 iovdd.n1352 iovdd.n120 0.0180786
R3808 iovdd.n1354 iovdd.n237 0.0180786
R3809 iovdd.n1356 iovdd.n114 0.0180786
R3810 iovdd.n1300 iovdd.n401 0.0180786
R3811 iovdd.n1298 iovdd.n400 0.0180786
R3812 iovdd.n1281 iovdd.n404 0.0180786
R3813 iovdd.n402 iovdd.n398 0.0180786
R3814 iovdd.n1280 iovdd.n407 0.0180786
R3815 iovdd.n405 iovdd.n396 0.0180786
R3816 iovdd.n1279 iovdd.n410 0.0180786
R3817 iovdd.n408 iovdd.n394 0.0180786
R3818 iovdd.n1303 iovdd.n1302 0.0180786
R3819 iovdd.n411 iovdd.n392 0.0180786
R3820 iovdd.n1305 iovdd.n390 0.0180786
R3821 iovdd.n1251 iovdd.n1249 0.0180786
R3822 iovdd.n1248 iovdd.n560 0.0180786
R3823 iovdd.n1254 iovdd.n1252 0.0180786
R3824 iovdd.n1246 iovdd.n561 0.0180786
R3825 iovdd.n1257 iovdd.n1255 0.0180786
R3826 iovdd.n1244 iovdd.n562 0.0180786
R3827 iovdd.n1260 iovdd.n1258 0.0180786
R3828 iovdd.n1242 iovdd.n563 0.0180786
R3829 iovdd.n1262 iovdd.n566 0.0180786
R3830 iovdd.n1263 iovdd.n565 0.0180786
R3831 iovdd.n564 iovdd.n388 0.0180786
R3832 iovdd.n786 iovdd.n785 0.0180786
R3833 iovdd.n784 iovdd.n775 0.0180786
R3834 iovdd.n788 iovdd.n787 0.0180786
R3835 iovdd.n783 iovdd.n776 0.0180786
R3836 iovdd.n1232 iovdd.n789 0.0180786
R3837 iovdd.n782 iovdd.n777 0.0180786
R3838 iovdd.n1234 iovdd.n779 0.0180786
R3839 iovdd.n1235 iovdd.n778 0.0180786
R3840 iovdd.n1237 iovdd.n569 0.0180786
R3841 iovdd.n773 iovdd.n568 0.0180786
R3842 iovdd.n770 iovdd.n387 0.0180786
R3843 iovdd.n399 iovdd.n56 0.0179603
R3844 iovdd.n227 iovdd.n69 0.0179603
R3845 iovdd.n197 iovdd.n90 0.0179603
R3846 iovdd.n176 iovdd.n103 0.0179603
R3847 iovdd.n1247 iovdd.n354 0.0179603
R3848 iovdd.n539 iovdd.n341 0.0179603
R3849 iovdd.n509 iovdd.n320 0.0179603
R3850 iovdd.n488 iovdd.n307 0.0179603
R3851 iovdd.n849 iovdd.n848 0.0179603
R3852 iovdd.n1175 iovdd.n833 0.0179603
R3853 iovdd.n1155 iovdd.n812 0.0179603
R3854 iovdd.n1141 iovdd.n799 0.0179603
R3855 iovdd.n1289 iovdd.n61 0.0175485
R3856 iovdd.n238 iovdd.n64 0.0175485
R3857 iovdd.n188 iovdd.n95 0.0175485
R3858 iovdd.n185 iovdd.n98 0.0175485
R3859 iovdd.n429 iovdd.n349 0.0175485
R3860 iovdd.n549 iovdd.n346 0.0175485
R3861 iovdd.n500 iovdd.n315 0.0175485
R3862 iovdd.n497 iovdd.n312 0.0175485
R3863 iovdd.n1191 iovdd.n841 0.0175485
R3864 iovdd.n1219 iovdd.n838 0.0175485
R3865 iovdd.n1149 iovdd.n807 0.0175485
R3866 iovdd.n1147 iovdd.n804 0.0175485
R3867 iovdd.n1311 iovdd.n296 0.0175485
R3868 iovdd.n133 iovdd.n78 0.0170873
R3869 iovdd.n135 iovdd.n81 0.0170873
R3870 iovdd.n447 iovdd.n332 0.0170873
R3871 iovdd.n449 iovdd.n329 0.0170873
R3872 iovdd.n1105 iovdd.n824 0.0170873
R3873 iovdd.n1107 iovdd.n821 0.0170873
R3874 iovdd.n403 iovdd.n55 0.0166755
R3875 iovdd.n125 iovdd.n70 0.0166755
R3876 iovdd.n143 iovdd.n89 0.0166755
R3877 iovdd.n159 iovdd.n104 0.0166755
R3878 iovdd.n1253 iovdd.n355 0.0166755
R3879 iovdd.n439 iovdd.n340 0.0166755
R3880 iovdd.n457 iovdd.n321 0.0166755
R3881 iovdd.n473 iovdd.n306 0.0166755
R3882 iovdd.n851 iovdd.n850 0.0166755
R3883 iovdd.n1097 iovdd.n832 0.0166755
R3884 iovdd.n1115 iovdd.n813 0.0166755
R3885 iovdd.n1131 iovdd.n798 0.0166755
R3886 iovdd.n397 iovdd.n53 0.0162143
R3887 iovdd.n224 iovdd.n72 0.0162143
R3888 iovdd.n200 iovdd.n87 0.0162143
R3889 iovdd.n173 iovdd.n106 0.0162143
R3890 iovdd.n1245 iovdd.n357 0.0162143
R3891 iovdd.n536 iovdd.n338 0.0162143
R3892 iovdd.n512 iovdd.n323 0.0162143
R3893 iovdd.n485 iovdd.n304 0.0162143
R3894 iovdd.n1230 iovdd.n791 0.0162143
R3895 iovdd.n1173 iovdd.n830 0.0162143
R3896 iovdd.n1157 iovdd.n815 0.0162143
R3897 iovdd.n1139 iovdd.n796 0.0162143
R3898 iovdd.n524 iovdd.n331 0.0158025
R3899 iovdd.n1165 iovdd.n822 0.0158025
R3900 iovdd.n212 iovdd.n79 0.0158025
R3901 iovdd.n235 iovdd.n62 0.0153413
R3902 iovdd.n235 iovdd.n63 0.0153413
R3903 iovdd.n151 iovdd.n96 0.0153413
R3904 iovdd.n151 iovdd.n97 0.0153413
R3905 iovdd.n432 iovdd.n348 0.0153413
R3906 iovdd.n432 iovdd.n347 0.0153413
R3907 iovdd.n465 iovdd.n314 0.0153413
R3908 iovdd.n465 iovdd.n313 0.0153413
R3909 iovdd.n1193 iovdd.n840 0.0153413
R3910 iovdd.n1193 iovdd.n839 0.0153413
R3911 iovdd.n1123 iovdd.n806 0.0153413
R3912 iovdd.n1123 iovdd.n805 0.0153413
R3913 iovdd.n1310 iovdd.n275 0.0153413
R3914 iovdd.n277 iovdd.n275 0.0153413
R3915 iovdd.n397 iovdd.n54 0.0144683
R3916 iovdd.n224 iovdd.n71 0.0144683
R3917 iovdd.n200 iovdd.n88 0.0144683
R3918 iovdd.n173 iovdd.n105 0.0144683
R3919 iovdd.n1245 iovdd.n356 0.0144683
R3920 iovdd.n536 iovdd.n339 0.0144683
R3921 iovdd.n512 iovdd.n322 0.0144683
R3922 iovdd.n485 iovdd.n305 0.0144683
R3923 iovdd.n852 iovdd.n791 0.0144683
R3924 iovdd.n1173 iovdd.n831 0.0144683
R3925 iovdd.n1157 iovdd.n814 0.0144683
R3926 iovdd.n1139 iovdd.n797 0.0144683
R3927 iovdd.n135 iovdd.n80 0.0135952
R3928 iovdd.n449 iovdd.n330 0.0135952
R3929 iovdd.n1105 iovdd.n823 0.0135952
R3930 iovdd.n116 iovdd 0.0127222
R3931 iovdd.n289 iovdd 0.0109762
R3932 iovdd.n1225 iovdd.n0 0.00923016
R3933 iovdd.n1228 iovdd.n1227 0.00835714
R3934 iovdd.n1357 iovdd.n45 0.00835714
R3935 iovdd.n1239 iovdd.n412 0.00748413
R3936 iovdd.n1357 iovdd.n112 0.00748413
R3937 iovdd.n1240 iovdd.n1239 0.00748413
R3938 iovdd.n298 iovdd.n275 0.00748413
R3939 iovdd.n1239 iovdd.n1238 0.00748413
R3940 iovdd.n1227 iovdd.n859 0.00748413
R3941 iovdd.n943 iovdd.n936 0.00740196
R3942 iovdd.n947 iovdd.n936 0.00740196
R3943 iovdd.n947 iovdd.n929 0.00740196
R3944 iovdd.n958 iovdd.n929 0.00740196
R3945 iovdd.n958 iovdd.n927 0.00740196
R3946 iovdd.n962 iovdd.n927 0.00740196
R3947 iovdd.n962 iovdd.n920 0.00740196
R3948 iovdd.n973 iovdd.n920 0.00740196
R3949 iovdd.n973 iovdd.n918 0.00740196
R3950 iovdd.n977 iovdd.n918 0.00740196
R3951 iovdd.n977 iovdd.n911 0.00740196
R3952 iovdd.n988 iovdd.n911 0.00740196
R3953 iovdd.n988 iovdd.n909 0.00740196
R3954 iovdd.n992 iovdd.n909 0.00740196
R3955 iovdd.n992 iovdd.n902 0.00740196
R3956 iovdd.n1003 iovdd.n902 0.00740196
R3957 iovdd.n1003 iovdd.n900 0.00740196
R3958 iovdd.n1007 iovdd.n900 0.00740196
R3959 iovdd.n1007 iovdd.n893 0.00740196
R3960 iovdd.n1018 iovdd.n893 0.00740196
R3961 iovdd.n1018 iovdd.n891 0.00740196
R3962 iovdd.n1022 iovdd.n891 0.00740196
R3963 iovdd.n1022 iovdd.n884 0.00740196
R3964 iovdd.n1033 iovdd.n884 0.00740196
R3965 iovdd.n1033 iovdd.n882 0.00740196
R3966 iovdd.n1037 iovdd.n882 0.00740196
R3967 iovdd.n1037 iovdd.n875 0.00740196
R3968 iovdd.n1048 iovdd.n875 0.00740196
R3969 iovdd.n1048 iovdd.n873 0.00740196
R3970 iovdd.n1052 iovdd.n873 0.00740196
R3971 iovdd.n1052 iovdd.n866 0.00740196
R3972 iovdd.n1063 iovdd.n866 0.00740196
R3973 iovdd.n1063 iovdd.n246 0.00740196
R3974 iovdd.n1315 iovdd.n246 0.00740196
R3975 iovdd.n1315 iovdd.n240 0.00740196
R3976 iovdd.n1327 iovdd.n240 0.00740196
R3977 iovdd.n1327 iovdd.n1326 0.00740196
R3978 iovdd.n946 iovdd.n945 0.00740196
R3979 iovdd.n946 iovdd.n928 0.00740196
R3980 iovdd.n959 iovdd.n928 0.00740196
R3981 iovdd.n960 iovdd.n959 0.00740196
R3982 iovdd.n961 iovdd.n960 0.00740196
R3983 iovdd.n961 iovdd.n919 0.00740196
R3984 iovdd.n974 iovdd.n919 0.00740196
R3985 iovdd.n975 iovdd.n974 0.00740196
R3986 iovdd.n976 iovdd.n975 0.00740196
R3987 iovdd.n976 iovdd.n910 0.00740196
R3988 iovdd.n989 iovdd.n910 0.00740196
R3989 iovdd.n990 iovdd.n989 0.00740196
R3990 iovdd.n991 iovdd.n990 0.00740196
R3991 iovdd.n991 iovdd.n901 0.00740196
R3992 iovdd.n1004 iovdd.n901 0.00740196
R3993 iovdd.n1005 iovdd.n1004 0.00740196
R3994 iovdd.n1006 iovdd.n1005 0.00740196
R3995 iovdd.n1006 iovdd.n892 0.00740196
R3996 iovdd.n1019 iovdd.n892 0.00740196
R3997 iovdd.n1020 iovdd.n1019 0.00740196
R3998 iovdd.n1021 iovdd.n1020 0.00740196
R3999 iovdd.n1021 iovdd.n883 0.00740196
R4000 iovdd.n1034 iovdd.n883 0.00740196
R4001 iovdd.n1035 iovdd.n1034 0.00740196
R4002 iovdd.n1036 iovdd.n1035 0.00740196
R4003 iovdd.n1036 iovdd.n874 0.00740196
R4004 iovdd.n1049 iovdd.n874 0.00740196
R4005 iovdd.n1050 iovdd.n1049 0.00740196
R4006 iovdd.n1051 iovdd.n1050 0.00740196
R4007 iovdd.n1051 iovdd.n865 0.00740196
R4008 iovdd.n1064 iovdd.n865 0.00740196
R4009 iovdd.n1314 iovdd.n247 0.00740196
R4010 iovdd.n1328 iovdd.n239 0.00740196
R4011 iovdd.n651 iovdd.n650 0.00740196
R4012 iovdd.n651 iovdd.n633 0.00740196
R4013 iovdd.n664 iovdd.n633 0.00740196
R4014 iovdd.n665 iovdd.n664 0.00740196
R4015 iovdd.n666 iovdd.n665 0.00740196
R4016 iovdd.n666 iovdd.n624 0.00740196
R4017 iovdd.n679 iovdd.n624 0.00740196
R4018 iovdd.n680 iovdd.n679 0.00740196
R4019 iovdd.n681 iovdd.n680 0.00740196
R4020 iovdd.n681 iovdd.n615 0.00740196
R4021 iovdd.n694 iovdd.n615 0.00740196
R4022 iovdd.n695 iovdd.n694 0.00740196
R4023 iovdd.n696 iovdd.n695 0.00740196
R4024 iovdd.n696 iovdd.n606 0.00740196
R4025 iovdd.n709 iovdd.n606 0.00740196
R4026 iovdd.n710 iovdd.n709 0.00740196
R4027 iovdd.n711 iovdd.n710 0.00740196
R4028 iovdd.n711 iovdd.n597 0.00740196
R4029 iovdd.n724 iovdd.n597 0.00740196
R4030 iovdd.n725 iovdd.n724 0.00740196
R4031 iovdd.n726 iovdd.n725 0.00740196
R4032 iovdd.n726 iovdd.n588 0.00740196
R4033 iovdd.n739 iovdd.n588 0.00740196
R4034 iovdd.n740 iovdd.n739 0.00740196
R4035 iovdd.n741 iovdd.n740 0.00740196
R4036 iovdd.n741 iovdd.n579 0.00740196
R4037 iovdd.n754 iovdd.n579 0.00740196
R4038 iovdd.n755 iovdd.n754 0.00740196
R4039 iovdd.n756 iovdd.n755 0.00740196
R4040 iovdd.n756 iovdd.n570 0.00740196
R4041 iovdd.n769 iovdd.n570 0.00740196
R4042 iovdd.n1265 iovdd.n422 0.00740196
R4043 iovdd.n1278 iovdd.n413 0.00740196
R4044 iovdd.n648 iovdd.n641 0.00740196
R4045 iovdd.n652 iovdd.n641 0.00740196
R4046 iovdd.n652 iovdd.n634 0.00740196
R4047 iovdd.n663 iovdd.n634 0.00740196
R4048 iovdd.n663 iovdd.n632 0.00740196
R4049 iovdd.n667 iovdd.n632 0.00740196
R4050 iovdd.n667 iovdd.n625 0.00740196
R4051 iovdd.n678 iovdd.n625 0.00740196
R4052 iovdd.n678 iovdd.n623 0.00740196
R4053 iovdd.n682 iovdd.n623 0.00740196
R4054 iovdd.n682 iovdd.n616 0.00740196
R4055 iovdd.n693 iovdd.n616 0.00740196
R4056 iovdd.n693 iovdd.n614 0.00740196
R4057 iovdd.n697 iovdd.n614 0.00740196
R4058 iovdd.n697 iovdd.n607 0.00740196
R4059 iovdd.n708 iovdd.n607 0.00740196
R4060 iovdd.n708 iovdd.n605 0.00740196
R4061 iovdd.n712 iovdd.n605 0.00740196
R4062 iovdd.n712 iovdd.n598 0.00740196
R4063 iovdd.n723 iovdd.n598 0.00740196
R4064 iovdd.n723 iovdd.n596 0.00740196
R4065 iovdd.n727 iovdd.n596 0.00740196
R4066 iovdd.n727 iovdd.n589 0.00740196
R4067 iovdd.n738 iovdd.n589 0.00740196
R4068 iovdd.n738 iovdd.n587 0.00740196
R4069 iovdd.n742 iovdd.n587 0.00740196
R4070 iovdd.n742 iovdd.n580 0.00740196
R4071 iovdd.n753 iovdd.n580 0.00740196
R4072 iovdd.n753 iovdd.n578 0.00740196
R4073 iovdd.n757 iovdd.n578 0.00740196
R4074 iovdd.n757 iovdd.n571 0.00740196
R4075 iovdd.n768 iovdd.n571 0.00740196
R4076 iovdd.n768 iovdd.n421 0.00740196
R4077 iovdd.n1266 iovdd.n421 0.00740196
R4078 iovdd.n1266 iovdd.n414 0.00740196
R4079 iovdd.n1277 iovdd.n414 0.00740196
R4080 iovdd.n1277 iovdd.n415 0.00740196
R4081 iovdd.n1355 iovdd 0.00671176
R4082 iovdd.n863 iovdd.n858 0.0057381
R4083 iovdd.n116 iovdd.n44 0.0057381
R4084 iovdd.n1353 iovdd.n1328 0.0047102
R4085 iovdd.n1301 iovdd.n1278 0.0047102
R4086 iovdd.n944 iovdd.n943 0.00442211
R4087 iovdd.n649 iovdd.n648 0.00442211
R4088 iovdd iovdd.n0 0.00399206
R4089 iovdd.n942 iovdd.n937 0.00395098
R4090 iovdd.n942 iovdd.n941 0.00395098
R4091 iovdd.n941 iovdd.n938 0.00395098
R4092 iovdd.n938 iovdd.n935 0.00395098
R4093 iovdd.n948 iovdd.n935 0.00395098
R4094 iovdd.n950 iovdd.n948 0.00395098
R4095 iovdd.n950 iovdd.n949 0.00395098
R4096 iovdd.n949 iovdd.n930 0.00395098
R4097 iovdd.n957 iovdd.n930 0.00395098
R4098 iovdd.n957 iovdd.n956 0.00395098
R4099 iovdd.n956 iovdd.n931 0.00395098
R4100 iovdd.n931 iovdd.n926 0.00395098
R4101 iovdd.n963 iovdd.n926 0.00395098
R4102 iovdd.n965 iovdd.n963 0.00395098
R4103 iovdd.n965 iovdd.n964 0.00395098
R4104 iovdd.n964 iovdd.n921 0.00395098
R4105 iovdd.n972 iovdd.n921 0.00395098
R4106 iovdd.n972 iovdd.n971 0.00395098
R4107 iovdd.n971 iovdd.n922 0.00395098
R4108 iovdd.n922 iovdd.n917 0.00395098
R4109 iovdd.n978 iovdd.n917 0.00395098
R4110 iovdd.n980 iovdd.n978 0.00395098
R4111 iovdd.n980 iovdd.n979 0.00395098
R4112 iovdd.n979 iovdd.n912 0.00395098
R4113 iovdd.n987 iovdd.n912 0.00395098
R4114 iovdd.n987 iovdd.n986 0.00395098
R4115 iovdd.n986 iovdd.n913 0.00395098
R4116 iovdd.n913 iovdd.n908 0.00395098
R4117 iovdd.n993 iovdd.n908 0.00395098
R4118 iovdd.n995 iovdd.n993 0.00395098
R4119 iovdd.n995 iovdd.n994 0.00395098
R4120 iovdd.n994 iovdd.n903 0.00395098
R4121 iovdd.n1002 iovdd.n903 0.00395098
R4122 iovdd.n1002 iovdd.n1001 0.00395098
R4123 iovdd.n1001 iovdd.n904 0.00395098
R4124 iovdd.n904 iovdd.n899 0.00395098
R4125 iovdd.n1008 iovdd.n899 0.00395098
R4126 iovdd.n1010 iovdd.n1008 0.00395098
R4127 iovdd.n1010 iovdd.n1009 0.00395098
R4128 iovdd.n1009 iovdd.n894 0.00395098
R4129 iovdd.n1017 iovdd.n894 0.00395098
R4130 iovdd.n1017 iovdd.n1016 0.00395098
R4131 iovdd.n1016 iovdd.n895 0.00395098
R4132 iovdd.n895 iovdd.n890 0.00395098
R4133 iovdd.n1023 iovdd.n890 0.00395098
R4134 iovdd.n1025 iovdd.n1023 0.00395098
R4135 iovdd.n1025 iovdd.n1024 0.00395098
R4136 iovdd.n1024 iovdd.n885 0.00395098
R4137 iovdd.n1032 iovdd.n885 0.00395098
R4138 iovdd.n1032 iovdd.n1031 0.00395098
R4139 iovdd.n1031 iovdd.n886 0.00395098
R4140 iovdd.n886 iovdd.n881 0.00395098
R4141 iovdd.n1038 iovdd.n881 0.00395098
R4142 iovdd.n1040 iovdd.n1038 0.00395098
R4143 iovdd.n1040 iovdd.n1039 0.00395098
R4144 iovdd.n1039 iovdd.n876 0.00395098
R4145 iovdd.n1047 iovdd.n876 0.00395098
R4146 iovdd.n1047 iovdd.n1046 0.00395098
R4147 iovdd.n1046 iovdd.n877 0.00395098
R4148 iovdd.n877 iovdd.n872 0.00395098
R4149 iovdd.n1053 iovdd.n872 0.00395098
R4150 iovdd.n1055 iovdd.n1053 0.00395098
R4151 iovdd.n1055 iovdd.n1054 0.00395098
R4152 iovdd.n1054 iovdd.n867 0.00395098
R4153 iovdd.n1062 iovdd.n867 0.00395098
R4154 iovdd.n1062 iovdd.n1061 0.00395098
R4155 iovdd.n1061 iovdd.n868 0.00395098
R4156 iovdd.n868 iovdd.n245 0.00395098
R4157 iovdd.n1316 iovdd.n245 0.00395098
R4158 iovdd.n1319 iovdd.n1316 0.00395098
R4159 iovdd.n1319 iovdd.n1318 0.00395098
R4160 iovdd.n1318 iovdd.n1317 0.00395098
R4161 iovdd.n1317 iovdd.n241 0.00395098
R4162 iovdd.n1325 iovdd.n241 0.00395098
R4163 iovdd.n647 iovdd.n642 0.00395098
R4164 iovdd.n647 iovdd.n646 0.00395098
R4165 iovdd.n646 iovdd.n643 0.00395098
R4166 iovdd.n643 iovdd.n640 0.00395098
R4167 iovdd.n653 iovdd.n640 0.00395098
R4168 iovdd.n655 iovdd.n653 0.00395098
R4169 iovdd.n655 iovdd.n654 0.00395098
R4170 iovdd.n654 iovdd.n635 0.00395098
R4171 iovdd.n662 iovdd.n635 0.00395098
R4172 iovdd.n662 iovdd.n661 0.00395098
R4173 iovdd.n661 iovdd.n636 0.00395098
R4174 iovdd.n636 iovdd.n631 0.00395098
R4175 iovdd.n668 iovdd.n631 0.00395098
R4176 iovdd.n670 iovdd.n668 0.00395098
R4177 iovdd.n670 iovdd.n669 0.00395098
R4178 iovdd.n669 iovdd.n626 0.00395098
R4179 iovdd.n677 iovdd.n626 0.00395098
R4180 iovdd.n677 iovdd.n676 0.00395098
R4181 iovdd.n676 iovdd.n627 0.00395098
R4182 iovdd.n627 iovdd.n622 0.00395098
R4183 iovdd.n683 iovdd.n622 0.00395098
R4184 iovdd.n685 iovdd.n683 0.00395098
R4185 iovdd.n685 iovdd.n684 0.00395098
R4186 iovdd.n684 iovdd.n617 0.00395098
R4187 iovdd.n692 iovdd.n617 0.00395098
R4188 iovdd.n692 iovdd.n691 0.00395098
R4189 iovdd.n691 iovdd.n618 0.00395098
R4190 iovdd.n618 iovdd.n613 0.00395098
R4191 iovdd.n698 iovdd.n613 0.00395098
R4192 iovdd.n700 iovdd.n698 0.00395098
R4193 iovdd.n700 iovdd.n699 0.00395098
R4194 iovdd.n699 iovdd.n608 0.00395098
R4195 iovdd.n707 iovdd.n608 0.00395098
R4196 iovdd.n707 iovdd.n706 0.00395098
R4197 iovdd.n706 iovdd.n609 0.00395098
R4198 iovdd.n609 iovdd.n604 0.00395098
R4199 iovdd.n713 iovdd.n604 0.00395098
R4200 iovdd.n715 iovdd.n713 0.00395098
R4201 iovdd.n715 iovdd.n714 0.00395098
R4202 iovdd.n714 iovdd.n599 0.00395098
R4203 iovdd.n722 iovdd.n599 0.00395098
R4204 iovdd.n722 iovdd.n721 0.00395098
R4205 iovdd.n721 iovdd.n600 0.00395098
R4206 iovdd.n600 iovdd.n595 0.00395098
R4207 iovdd.n728 iovdd.n595 0.00395098
R4208 iovdd.n730 iovdd.n728 0.00395098
R4209 iovdd.n730 iovdd.n729 0.00395098
R4210 iovdd.n729 iovdd.n590 0.00395098
R4211 iovdd.n737 iovdd.n590 0.00395098
R4212 iovdd.n737 iovdd.n736 0.00395098
R4213 iovdd.n736 iovdd.n591 0.00395098
R4214 iovdd.n591 iovdd.n586 0.00395098
R4215 iovdd.n743 iovdd.n586 0.00395098
R4216 iovdd.n745 iovdd.n743 0.00395098
R4217 iovdd.n745 iovdd.n744 0.00395098
R4218 iovdd.n744 iovdd.n581 0.00395098
R4219 iovdd.n752 iovdd.n581 0.00395098
R4220 iovdd.n752 iovdd.n751 0.00395098
R4221 iovdd.n751 iovdd.n582 0.00395098
R4222 iovdd.n582 iovdd.n577 0.00395098
R4223 iovdd.n758 iovdd.n577 0.00395098
R4224 iovdd.n760 iovdd.n758 0.00395098
R4225 iovdd.n760 iovdd.n759 0.00395098
R4226 iovdd.n759 iovdd.n572 0.00395098
R4227 iovdd.n767 iovdd.n572 0.00395098
R4228 iovdd.n767 iovdd.n766 0.00395098
R4229 iovdd.n766 iovdd.n573 0.00395098
R4230 iovdd.n573 iovdd.n420 0.00395098
R4231 iovdd.n1267 iovdd.n420 0.00395098
R4232 iovdd.n1269 iovdd.n1267 0.00395098
R4233 iovdd.n1269 iovdd.n1268 0.00395098
R4234 iovdd.n1268 iovdd.n416 0.00395098
R4235 iovdd.n1276 iovdd.n416 0.00395098
R4236 iovdd.n1276 iovdd.n1275 0.00395098
R4237 iovdd.n1239 iovdd.n49 0.00360916
R4238 iovdd.n1306 iovdd.n375 0.00339474
R4239 iovdd.n1218 iovdd.n247 0.00326078
R4240 iovdd.n1233 iovdd.n422 0.00326078
R4241 iovdd.n1314 iovdd.n1313 0.00298471
R4242 iovdd.n1265 iovdd.n1264 0.00298471
R4243 iovdd.n772 iovdd.n375 0.00285867
R4244 iovdd.n1274 iovdd 0.00261765
R4245 iovdd.n290 iovdd.n289 0.00224603
R4246 iovdd.n1236 iovdd.n774 0.00219098
R4247 iovdd.n1264 iovdd.n559 0.00219098
R4248 iovdd.n1261 iovdd.n559 0.00219098
R4249 iovdd.n1273 iovdd 0.00196667
R4250 iovdd.n1323 iovdd 0.00196667
R4251 iovdd.n940 iovdd.n934 0.00191176
R4252 iovdd.n951 iovdd.n934 0.00191176
R4253 iovdd.n951 iovdd.n932 0.00191176
R4254 iovdd.n955 iovdd.n932 0.00191176
R4255 iovdd.n955 iovdd.n925 0.00191176
R4256 iovdd.n966 iovdd.n925 0.00191176
R4257 iovdd.n966 iovdd.n923 0.00191176
R4258 iovdd.n970 iovdd.n923 0.00191176
R4259 iovdd.n970 iovdd.n916 0.00191176
R4260 iovdd.n981 iovdd.n916 0.00191176
R4261 iovdd.n981 iovdd.n914 0.00191176
R4262 iovdd.n985 iovdd.n914 0.00191176
R4263 iovdd.n985 iovdd.n907 0.00191176
R4264 iovdd.n996 iovdd.n907 0.00191176
R4265 iovdd.n996 iovdd.n905 0.00191176
R4266 iovdd.n1000 iovdd.n905 0.00191176
R4267 iovdd.n1000 iovdd.n898 0.00191176
R4268 iovdd.n1011 iovdd.n898 0.00191176
R4269 iovdd.n1011 iovdd.n896 0.00191176
R4270 iovdd.n1015 iovdd.n896 0.00191176
R4271 iovdd.n1015 iovdd.n889 0.00191176
R4272 iovdd.n1026 iovdd.n889 0.00191176
R4273 iovdd.n1026 iovdd.n887 0.00191176
R4274 iovdd.n1030 iovdd.n887 0.00191176
R4275 iovdd.n1030 iovdd.n880 0.00191176
R4276 iovdd.n1041 iovdd.n880 0.00191176
R4277 iovdd.n1041 iovdd.n878 0.00191176
R4278 iovdd.n1045 iovdd.n878 0.00191176
R4279 iovdd.n1045 iovdd.n871 0.00191176
R4280 iovdd.n1056 iovdd.n871 0.00191176
R4281 iovdd.n1056 iovdd.n869 0.00191176
R4282 iovdd.n1060 iovdd.n869 0.00191176
R4283 iovdd.n1060 iovdd.n244 0.00191176
R4284 iovdd.n1320 iovdd.n244 0.00191176
R4285 iovdd.n1320 iovdd.n242 0.00191176
R4286 iovdd.n1324 iovdd.n242 0.00191176
R4287 iovdd.n645 iovdd.n639 0.00191176
R4288 iovdd.n656 iovdd.n639 0.00191176
R4289 iovdd.n656 iovdd.n637 0.00191176
R4290 iovdd.n660 iovdd.n637 0.00191176
R4291 iovdd.n660 iovdd.n630 0.00191176
R4292 iovdd.n671 iovdd.n630 0.00191176
R4293 iovdd.n671 iovdd.n628 0.00191176
R4294 iovdd.n675 iovdd.n628 0.00191176
R4295 iovdd.n675 iovdd.n621 0.00191176
R4296 iovdd.n686 iovdd.n621 0.00191176
R4297 iovdd.n686 iovdd.n619 0.00191176
R4298 iovdd.n690 iovdd.n619 0.00191176
R4299 iovdd.n690 iovdd.n612 0.00191176
R4300 iovdd.n701 iovdd.n612 0.00191176
R4301 iovdd.n701 iovdd.n610 0.00191176
R4302 iovdd.n705 iovdd.n610 0.00191176
R4303 iovdd.n705 iovdd.n603 0.00191176
R4304 iovdd.n716 iovdd.n603 0.00191176
R4305 iovdd.n716 iovdd.n601 0.00191176
R4306 iovdd.n720 iovdd.n601 0.00191176
R4307 iovdd.n720 iovdd.n594 0.00191176
R4308 iovdd.n731 iovdd.n594 0.00191176
R4309 iovdd.n731 iovdd.n592 0.00191176
R4310 iovdd.n735 iovdd.n592 0.00191176
R4311 iovdd.n735 iovdd.n585 0.00191176
R4312 iovdd.n746 iovdd.n585 0.00191176
R4313 iovdd.n746 iovdd.n583 0.00191176
R4314 iovdd.n750 iovdd.n583 0.00191176
R4315 iovdd.n750 iovdd.n576 0.00191176
R4316 iovdd.n761 iovdd.n576 0.00191176
R4317 iovdd.n761 iovdd.n574 0.00191176
R4318 iovdd.n765 iovdd.n574 0.00191176
R4319 iovdd.n765 iovdd.n419 0.00191176
R4320 iovdd.n1270 iovdd.n419 0.00191176
R4321 iovdd.n1270 iovdd.n417 0.00191176
R4322 iovdd.n1274 iovdd.n417 0.00191176
R4323 iovdd.n1294 iovdd.n389 0.00189683
R4324 iovdd.n1286 iovdd.n115 0.00189683
R4325 iovdd.n1183 iovdd.n774 0.00189683
R4326 iovdd.n1221 iovdd.n1090 0.00189683
R4327 iovdd.n559 iovdd.n558 0.00189683
R4328 iovdd.n552 iovdd.n431 0.00189683
R4329 iovdd.n1222 iovdd.n1221 0.00184541
R4330 iovdd.n1218 iovdd.n864 0.00184541
R4331 iovdd.n431 iovdd.n248 0.00184541
R4332 iovdd.n548 iovdd.n431 0.00184541
R4333 iovdd.n1329 iovdd.n115 0.00184541
R4334 iovdd.n548 iovdd.n547 0.00184541
R4335 iovdd.n1313 iovdd.n248 0.00184541
R4336 iovdd.n1223 iovdd.n1222 0.00184541
R4337 iovdd.n1221 iovdd.n864 0.00184541
R4338 iovdd.n1353 iovdd.n1329 0.00184541
R4339 iovdd.n1233 iovdd.n781 0.00184541
R4340 iovdd.n1297 iovdd.n389 0.00184541
R4341 iovdd.n1301 iovdd.n1297 0.00184541
R4342 iovdd.n781 iovdd.n774 0.00184541
R4343 iovdd.n772 iovdd.n49 0.00178655
R4344 iovdd.n940 iovdd.n939 0.0016983
R4345 iovdd.n645 iovdd.n644 0.0016983
R4346 iovdd.n547 iovdd.n239 0.00153529
R4347 iovdd.n1261 iovdd.n413 0.00153529
R4348 iovdd.n118 iovdd.n115 0.00150078
R4349 iovdd.n391 iovdd.n389 0.00150078
R4350 iovdd.n657 iovdd.n638 0.00147778
R4351 iovdd.n658 iovdd.n657 0.00147778
R4352 iovdd.n659 iovdd.n658 0.00147778
R4353 iovdd.n659 iovdd.n629 0.00147778
R4354 iovdd.n672 iovdd.n629 0.00147778
R4355 iovdd.n673 iovdd.n672 0.00147778
R4356 iovdd.n674 iovdd.n673 0.00147778
R4357 iovdd.n674 iovdd.n620 0.00147778
R4358 iovdd.n687 iovdd.n620 0.00147778
R4359 iovdd.n688 iovdd.n687 0.00147778
R4360 iovdd.n689 iovdd.n688 0.00147778
R4361 iovdd.n689 iovdd.n611 0.00147778
R4362 iovdd.n702 iovdd.n611 0.00147778
R4363 iovdd.n703 iovdd.n702 0.00147778
R4364 iovdd.n704 iovdd.n703 0.00147778
R4365 iovdd.n704 iovdd.n602 0.00147778
R4366 iovdd.n717 iovdd.n602 0.00147778
R4367 iovdd.n718 iovdd.n717 0.00147778
R4368 iovdd.n719 iovdd.n718 0.00147778
R4369 iovdd.n719 iovdd.n593 0.00147778
R4370 iovdd.n732 iovdd.n593 0.00147778
R4371 iovdd.n733 iovdd.n732 0.00147778
R4372 iovdd.n734 iovdd.n733 0.00147778
R4373 iovdd.n734 iovdd.n584 0.00147778
R4374 iovdd.n747 iovdd.n584 0.00147778
R4375 iovdd.n748 iovdd.n747 0.00147778
R4376 iovdd.n749 iovdd.n748 0.00147778
R4377 iovdd.n749 iovdd.n575 0.00147778
R4378 iovdd.n762 iovdd.n575 0.00147778
R4379 iovdd.n763 iovdd.n762 0.00147778
R4380 iovdd.n764 iovdd.n763 0.00147778
R4381 iovdd.n764 iovdd.n418 0.00147778
R4382 iovdd.n1271 iovdd.n418 0.00147778
R4383 iovdd.n1272 iovdd.n1271 0.00147778
R4384 iovdd.n1273 iovdd.n1272 0.00147778
R4385 iovdd.n952 iovdd.n933 0.00147778
R4386 iovdd.n953 iovdd.n952 0.00147778
R4387 iovdd.n954 iovdd.n953 0.00147778
R4388 iovdd.n954 iovdd.n924 0.00147778
R4389 iovdd.n967 iovdd.n924 0.00147778
R4390 iovdd.n968 iovdd.n967 0.00147778
R4391 iovdd.n969 iovdd.n968 0.00147778
R4392 iovdd.n969 iovdd.n915 0.00147778
R4393 iovdd.n982 iovdd.n915 0.00147778
R4394 iovdd.n983 iovdd.n982 0.00147778
R4395 iovdd.n984 iovdd.n983 0.00147778
R4396 iovdd.n984 iovdd.n906 0.00147778
R4397 iovdd.n997 iovdd.n906 0.00147778
R4398 iovdd.n998 iovdd.n997 0.00147778
R4399 iovdd.n999 iovdd.n998 0.00147778
R4400 iovdd.n999 iovdd.n897 0.00147778
R4401 iovdd.n1012 iovdd.n897 0.00147778
R4402 iovdd.n1013 iovdd.n1012 0.00147778
R4403 iovdd.n1014 iovdd.n1013 0.00147778
R4404 iovdd.n1014 iovdd.n888 0.00147778
R4405 iovdd.n1027 iovdd.n888 0.00147778
R4406 iovdd.n1028 iovdd.n1027 0.00147778
R4407 iovdd.n1029 iovdd.n1028 0.00147778
R4408 iovdd.n1029 iovdd.n879 0.00147778
R4409 iovdd.n1042 iovdd.n879 0.00147778
R4410 iovdd.n1043 iovdd.n1042 0.00147778
R4411 iovdd.n1044 iovdd.n1043 0.00147778
R4412 iovdd.n1044 iovdd.n870 0.00147778
R4413 iovdd.n1057 iovdd.n870 0.00147778
R4414 iovdd.n1058 iovdd.n1057 0.00147778
R4415 iovdd.n1059 iovdd.n1058 0.00147778
R4416 iovdd.n1059 iovdd.n243 0.00147778
R4417 iovdd.n1321 iovdd.n243 0.00147778
R4418 iovdd.n1322 iovdd.n1321 0.00147778
R4419 iovdd.n1323 iovdd.n1322 0.00147778
R4420 iovdd.n1223 iovdd.n1064 0.00125922
R4421 iovdd.n1236 iovdd.n769 0.00125922
R4422 iovdd.n1307 iovdd.n1306 0.00125049
R4423 iovdd.n1355 iovdd.n118 0.0011902
R4424 iovdd.n1304 iovdd.n391 0.0011902
R4425 iovdd.n1360 iovdd.n1359 0.00101087
R4426 iovdd.n1309 iovdd.n25 0.001
R4427 iovdd.n1229 iovdd.n8 0.001
R4428 iovdd.n363 iovdd.n7 0.001
R4429 iovdd.n376 iovdd.n7 0.001
R4430 iovdd.n857 iovdd.n9 0.001
R4431 iovdd.n377 iovdd.n9 0.001
R4432 iovdd.n364 iovdd.n11 0.001
R4433 iovdd.n378 iovdd.n11 0.001
R4434 iovdd.n365 iovdd.n13 0.001
R4435 iovdd.n379 iovdd.n13 0.001
R4436 iovdd.n366 iovdd.n17 0.001
R4437 iovdd.n380 iovdd.n17 0.001
R4438 iovdd.n367 iovdd.n20 0.001
R4439 iovdd.n381 iovdd.n20 0.001
R4440 iovdd.n368 iovdd.n23 0.001
R4441 iovdd.n1308 iovdd.n23 0.001
R4442 iovdd.n1309 iovdd.n362 0.001
R4443 iovdd.n369 iovdd.n28 0.001
R4444 iovdd.n382 iovdd.n28 0.001
R4445 iovdd.n370 iovdd.n31 0.001
R4446 iovdd.n383 iovdd.n31 0.001
R4447 iovdd.n371 iovdd.n34 0.001
R4448 iovdd.n384 iovdd.n34 0.001
R4449 iovdd.n372 iovdd.n37 0.001
R4450 iovdd.n385 iovdd.n37 0.001
R4451 iovdd.n373 iovdd.n40 0.001
R4452 iovdd.n386 iovdd.n40 0.001
R4453 iovdd.n1359 iovdd.n48 0.001
R4454 iovdd.n1359 iovdd.n47 0.001
R4455 iovdd.n374 iovdd.n43 0.001
R4456 iovdd.n47 iovdd.n4 0.001
R4457 iovdd.n386 iovdd.n42 0.001
R4458 iovdd.n385 iovdd.n39 0.001
R4459 iovdd.n384 iovdd.n36 0.001
R4460 iovdd.n383 iovdd.n33 0.001
R4461 iovdd.n382 iovdd.n30 0.001
R4462 iovdd.n362 iovdd.n27 0.001
R4463 iovdd.n1309 iovdd.n1308 0.001
R4464 iovdd.n381 iovdd.n22 0.001
R4465 iovdd.n380 iovdd.n19 0.001
R4466 iovdd.n379 iovdd.n16 0.001
R4467 iovdd.n378 iovdd.n12 0.001
R4468 iovdd.n377 iovdd.n10 0.001
R4469 iovdd.n1229 iovdd.n376 0.001
R4470 iovdd.n374 iovdd.n4 0.001
R4471 iovdd.n48 iovdd.n42 0.001
R4472 iovdd.n373 iovdd.n39 0.001
R4473 iovdd.n372 iovdd.n36 0.001
R4474 iovdd.n371 iovdd.n33 0.001
R4475 iovdd.n370 iovdd.n30 0.001
R4476 iovdd.n369 iovdd.n27 0.001
R4477 iovdd.n368 iovdd.n22 0.001
R4478 iovdd.n367 iovdd.n19 0.001
R4479 iovdd.n366 iovdd.n16 0.001
R4480 iovdd.n365 iovdd.n12 0.001
R4481 iovdd.n364 iovdd.n10 0.001
R4482 iovdd.n1229 iovdd.n857 0.001
R4483 iovdd.n363 iovdd.n5 0.001
R4484 iovdd.n8 iovdd.n3 0.001
R4485 iovdd.n1361 iovdd.n3 0.001
R4486 iovdd.n1362 iovdd.n2 0.001
R4487 iovdd.n15 iovdd.n14 0.001
R4488 iovdd.n293 iovdd.n18 0.001
R4489 iovdd.n292 iovdd.n21 0.001
R4490 iovdd.n291 iovdd.n24 0.001
R4491 iovdd.n288 iovdd.n25 0.001
R4492 iovdd.n288 iovdd.n26 0.001
R4493 iovdd.n286 iovdd.n29 0.001
R4494 iovdd.n284 iovdd.n32 0.001
R4495 iovdd.n282 iovdd.n35 0.001
R4496 iovdd.n280 iovdd.n38 0.001
R4497 iovdd.n278 iovdd.n41 0.001
R4498 iovdd.n1359 iovdd.n41 0.001
R4499 iovdd.n278 iovdd.n38 0.001
R4500 iovdd.n280 iovdd.n35 0.001
R4501 iovdd.n282 iovdd.n32 0.001
R4502 iovdd.n284 iovdd.n29 0.001
R4503 iovdd.n286 iovdd.n26 0.001
R4504 iovdd.n1309 iovdd.n24 0.001
R4505 iovdd.n1229 iovdd.n6 0.001
R4506 iovdd.n291 iovdd.n21 0.001
R4507 iovdd.n292 iovdd.n18 0.001
R4508 iovdd.n293 iovdd.n15 0.001
R4509 iovdd.n14 iovdd.n2 0.001
R4510 iovdd.n1362 iovdd.n1361 0.001
R4511 vdd.n74 vdd.n73 1.50539
R4512 vdd.n1 vdd.n0 1.5005
R4513 vdd.n69 vdd.n68 1.5005
R4514 vdd.n67 vdd.n66 1.5005
R4515 vdd.n5 vdd.n4 1.5005
R4516 vdd.n61 vdd.n60 1.5005
R4517 vdd.n59 vdd.n58 1.5005
R4518 vdd.n9 vdd.n8 1.5005
R4519 vdd.n53 vdd.n52 1.5005
R4520 vdd.n51 vdd.n50 1.5005
R4521 vdd.n13 vdd.n12 1.5005
R4522 vdd.n45 vdd.n44 1.5005
R4523 vdd.n43 vdd.n42 1.5005
R4524 vdd.n17 vdd.n16 1.5005
R4525 vdd.n37 vdd.n36 1.5005
R4526 vdd.n35 vdd.n34 1.5005
R4527 vdd.n21 vdd.n20 1.5005
R4528 vdd.n29 vdd.n28 1.5005
R4529 vdd.n27 vdd.n26 1.5005
R4530 vdd.n75 vdd 0.6957
R4531 vdd.n73 vdd.n72 0.314786
R4532 vdd.n71 vdd.n70 0.314786
R4533 vdd.n3 vdd.n2 0.314786
R4534 vdd.n65 vdd.n64 0.314786
R4535 vdd.n63 vdd.n62 0.314786
R4536 vdd.n7 vdd.n6 0.314786
R4537 vdd.n57 vdd.n56 0.314786
R4538 vdd.n55 vdd.n54 0.314786
R4539 vdd.n11 vdd.n10 0.314786
R4540 vdd.n49 vdd.n48 0.314786
R4541 vdd.n47 vdd.n46 0.314786
R4542 vdd.n15 vdd.n14 0.314786
R4543 vdd.n41 vdd.n40 0.314786
R4544 vdd.n39 vdd.n38 0.314786
R4545 vdd.n19 vdd.n18 0.314786
R4546 vdd.n33 vdd.n32 0.314786
R4547 vdd.n31 vdd.n30 0.314786
R4548 vdd.n23 vdd.n22 0.314786
R4549 vdd.n24 vdd 0.217715
R4550 vdd.n51 vdd 0.195018
R4551 vdd.n25 vdd.n24 0.146103
R4552 vdd.n26 vdd.n25 0.0354467
R4553 vdd.n25 vdd.n22 0.0314255
R4554 vdd.n28 vdd.n27 0.00921287
R4555 vdd.n28 vdd.n20 0.00921287
R4556 vdd.n35 vdd.n20 0.00921287
R4557 vdd.n36 vdd.n35 0.00921287
R4558 vdd.n36 vdd.n16 0.00921287
R4559 vdd.n43 vdd.n16 0.00921287
R4560 vdd.n44 vdd.n43 0.00921287
R4561 vdd.n44 vdd.n12 0.00921287
R4562 vdd.n51 vdd.n12 0.00921287
R4563 vdd.n52 vdd.n51 0.00921287
R4564 vdd.n52 vdd.n8 0.00921287
R4565 vdd.n59 vdd.n8 0.00921287
R4566 vdd.n60 vdd.n59 0.00921287
R4567 vdd.n60 vdd.n4 0.00921287
R4568 vdd.n67 vdd.n4 0.00921287
R4569 vdd.n68 vdd.n67 0.00921287
R4570 vdd.n68 vdd.n0 0.00921287
R4571 vdd.n74 vdd.n0 0.00921287
R4572 vdd.n26 vdd.n23 0.00538889
R4573 vdd.n29 vdd.n23 0.00538889
R4574 vdd.n30 vdd.n29 0.00538889
R4575 vdd.n30 vdd.n21 0.00538889
R4576 vdd.n33 vdd.n21 0.00538889
R4577 vdd.n34 vdd.n33 0.00538889
R4578 vdd.n34 vdd.n19 0.00538889
R4579 vdd.n37 vdd.n19 0.00538889
R4580 vdd.n38 vdd.n37 0.00538889
R4581 vdd.n38 vdd.n17 0.00538889
R4582 vdd.n41 vdd.n17 0.00538889
R4583 vdd.n42 vdd.n41 0.00538889
R4584 vdd.n42 vdd.n15 0.00538889
R4585 vdd.n45 vdd.n15 0.00538889
R4586 vdd.n46 vdd.n45 0.00538889
R4587 vdd.n46 vdd.n13 0.00538889
R4588 vdd.n49 vdd.n13 0.00538889
R4589 vdd.n50 vdd.n49 0.00538889
R4590 vdd.n50 vdd.n11 0.00538889
R4591 vdd.n53 vdd.n11 0.00538889
R4592 vdd.n54 vdd.n53 0.00538889
R4593 vdd.n54 vdd.n9 0.00538889
R4594 vdd.n57 vdd.n9 0.00538889
R4595 vdd.n58 vdd.n57 0.00538889
R4596 vdd.n58 vdd.n7 0.00538889
R4597 vdd.n61 vdd.n7 0.00538889
R4598 vdd.n62 vdd.n61 0.00538889
R4599 vdd.n62 vdd.n5 0.00538889
R4600 vdd.n65 vdd.n5 0.00538889
R4601 vdd.n66 vdd.n65 0.00538889
R4602 vdd.n66 vdd.n3 0.00538889
R4603 vdd.n69 vdd.n3 0.00538889
R4604 vdd.n70 vdd.n69 0.00538889
R4605 vdd.n70 vdd.n1 0.00538889
R4606 vdd.n73 vdd.n1 0.00538889
R4607 vdd.n27 vdd.n24 0.00485644
R4608 vdd.n75 vdd.n74 0.00485644
R4609 vdd vdd.n75 0.00485644
R4610 vdd.n72 vdd 0.0035
R4611 vdd.n31 vdd.n22 0.0025
R4612 vdd.n32 vdd.n31 0.0025
R4613 vdd.n32 vdd.n18 0.0025
R4614 vdd.n39 vdd.n18 0.0025
R4615 vdd.n40 vdd.n39 0.0025
R4616 vdd.n40 vdd.n14 0.0025
R4617 vdd.n47 vdd.n14 0.0025
R4618 vdd.n48 vdd.n47 0.0025
R4619 vdd.n48 vdd.n10 0.0025
R4620 vdd.n55 vdd.n10 0.0025
R4621 vdd.n56 vdd.n55 0.0025
R4622 vdd.n56 vdd.n6 0.0025
R4623 vdd.n63 vdd.n6 0.0025
R4624 vdd.n64 vdd.n63 0.0025
R4625 vdd.n64 vdd.n2 0.0025
R4626 vdd.n71 vdd.n2 0.0025
R4627 vdd.n72 vdd.n71 0.0025
C0 sg13g2_DCNDiode_0.guard iovdd 0.1269f
C1 iovdd iovss 0.31233p
C2 vdd iovss 0.24767p
C3 sg13g2_DCNDiode_0.guard iovss 0.26938p $ **FLOATING
.ends

