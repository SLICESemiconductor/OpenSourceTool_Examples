* Extracted by KLayout with SG13G2 LVS runset on : 29/08/2025 17:54

.SUBCKT OTA_final vssa vtail vinn vout vinp pdio vdda
M$1 vssa vssa vssa vssa sg13_lv_nmos L=1u W=8u AS=2.2p AD=2.12p PS=16.4u
+ PD=16.24u
M$2 vssa vssa vssa vssa sg13_lv_nmos L=2u W=12u AS=2.28p AD=2.28p PS=16.56u
+ PD=16.56u
M$4 vssa vssa \$49 vssa sg13_lv_nmos L=2u W=2u AS=0.38p AD=0.38p PS=2.76u
+ PD=2.76u
M$12 vssa \$13 vtail vssa sg13_lv_nmos L=2u W=8u AS=1.52p AD=1.52p PS=11.04u
+ PD=11.04u
M$14 vssa \$13 \$13 vssa sg13_lv_nmos L=2u W=8u AS=1.52p AD=1.52p PS=11.04u
+ PD=11.04u
M$34 vssa vssa \$10 vssa sg13_lv_nmos L=2u W=2u AS=0.38p AD=0.38p PS=2.76u
+ PD=2.76u
M$41 vdda vdda vdda vdda sg13_lv_pmos L=1u W=8u AS=2.12p AD=2.12p PS=16.24u
+ PD=16.24u
M$42 vdda vdda vdda vdda sg13_lv_pmos L=2u W=16u AS=3.04p AD=3.04p PS=22.08u
+ PD=22.08u
M$52 vdda pdio vout vdda sg13_lv_pmos L=2u W=8u AS=1.52p AD=1.52p PS=11.04u
+ PD=11.04u
M$54 vdda pdio pdio vdda sg13_lv_pmos L=2u W=8u AS=1.52p AD=1.52p PS=11.04u
+ PD=11.04u
M$81 vtail vtail vtail vtail sg13_lv_nmos L=0.5u W=32u AS=6.38p AD=6.38p
+ PS=46.76u PD=46.76u
M$113 vtail vinp pdio vtail sg13_lv_nmos L=0.5u W=32u AS=6.38p AD=6.38p
+ PS=46.76u PD=46.76u
M$121 vtail vinn vout vtail sg13_lv_nmos L=0.5u W=32u AS=6.38p AD=6.38p
+ PS=46.76u PD=46.76u
.ENDS OTA_final
