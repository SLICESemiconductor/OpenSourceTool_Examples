** sch_path: /usr/local/share/xschem/xschem_library/devices/loopgainprobe.sch
**.subckt loopgainprobe a b
*.iopin b
*.iopin a
**** begin user architecture code

Ii

Ii 0 x DC 0 AC 0
Vi x a DC 0 AC 1
Vnodebuffer b x 0
**** end user architecture code
**.ends
.end
