* NGSPICE file created from sg13g2_IOPadTriOut30mA_flat.ext - technology: ihp-sg13g2

.subckt sg13g2_IOPadTriOut30mA_flat c2p_en c2p pad vdd vss iovdd iovss
X0 sg13g2_GateDecode_0.pgate.t2 iovdd.t0 dpantenna l=0.78u w=0.78u
X1 iovdd.t14 sg13g2_GateDecode_0.pgate.t3 pad.t10 iovdd.t0 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X2 iovdd.t11 sg13g2_GateDecode_0.pgate.t4 pad.t13 iovdd.t0 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X3 iovss sg13g2_GateDecode_0.ngate.t2 pad.t21 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X4 pad.t5 sg13g2_GateDecode_0.pgate.t5 iovdd.t28 iovdd.t0 sg13_hv_pmos ad=3.9294p pd=7.84u as=3.1302p ps=14.26u w=6.66u l=0.6u
X5 iovdd.t8 sg13g2_GateDecode_0.pgate.t6 pad.t8 iovdd.t0 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X6 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t1 c2p_en.t0 a_8230_33842# iovss sg13_lv_nmos ad=1.4148p pd=8.58u as=0.7467p ps=4.31u w=3.93u l=0.13u
X7 pad.t15 sg13g2_GateDecode_0.pgate.t7 iovdd.t16 iovdd.t0 sg13_hv_pmos ad=4.9284p pd=14.8u as=2.1312p ps=7.3u w=6.66u l=0.6u
X8 iovdd.t15 sg13g2_GateDecode_0.pgate.t4 pad.t12 iovdd.t0 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X9 iovss pad.t24 dantenna l=1.26u w=27.78u
X10 pad.t23 sg13g2_GateDecode_0.ngate.t3 iovss iovss sg13_hv_nmos ad=3.256p pd=10.28u as=1.408p ps=5.04u w=4.4u l=0.6u
X11 pad.t17 sg13g2_GateDecode_0.ngate.t4 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X12 iovss sg13g2_GateDecode_0.ngate.t5 pad.t18 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X13 iovss sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq iovss sg13_lv_nmos ad=1.4148p pd=8.58u as=0.7467p ps=4.31u w=3.93u l=0.13u
X14 a_7724_30170# sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq iovss iovss sg13_hv_nmos ad=0.646p pd=4.48u as=0.361p ps=2.28u w=1.9u l=0.45u
X15 iovdd a_7724_30170# a_7656_30206# iovdd sg13_hv_pmos ad=57f pd=0.68u as=0.102p ps=1.28u w=0.3u l=0.45u
X16 pad.t4 sg13g2_GateDecode_0.pgate.t5 iovdd.t25 iovdd.t0 sg13_hv_pmos ad=3.9294p pd=7.84u as=3.1302p ps=14.26u w=6.66u l=0.6u
X17 iovdd.t1 sg13g2_GateDecode_0.pgate.t6 pad.t7 iovdd.t0 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X18 iovdd.t5 sg13g2_GateDecode_0.pgate.t8 pad.t11 iovdd.t0 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X19 iovss sg13g2_GateDecode_0.ngate.t6 pad.t22 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X20 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t0 c2p.t0 vdd.t8 vdd.t2 sg13_lv_pmos ad=0.8379p pd=4.79u as=1.4994p ps=9.5u w=4.41u l=0.13u
X21 sg13g2_GateDecode_0.ngate.t0 a_7724_30170# iovdd iovdd sg13_hv_pmos ad=1.326p pd=8.48u as=1.326p ps=8.48u w=3.9u l=0.45u
X22 pad.t14 sg13g2_GateDecode_0.pgate.t7 iovdd.t13 iovdd.t0 sg13_hv_pmos ad=4.9284p pd=14.8u as=2.1312p ps=7.3u w=6.66u l=0.6u
X23 iovdd.t12 sg13g2_GateDecode_0.pgate.t9 pad.t2 iovdd.t0 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X24 a_8426_30170# a_8358_30206# iovdd iovdd sg13_hv_pmos ad=0.102p pd=1.28u as=57f ps=0.68u w=0.3u l=0.45u
X25 a_7750_34876# c2p.t1 vdd.t7 vdd.t4 sg13_lv_pmos ad=0.8379p pd=4.79u as=1.4994p ps=9.5u w=4.41u l=0.13u
X26 iovdd.t6 sg13g2_GateDecode_0.pgate.t8 pad.t9 iovdd.t0 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X27 pad.t13 sg13g2_GateDecode_0.pgate.t10 iovdd.t7 iovdd.t0 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X28 pad.t19 sg13g2_GateDecode_0.ngate.t7 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X29 iovss sg13g2_GateDecode_0.ngate.t8 pad.t16 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X30 pad.t18 sg13g2_GateDecode_0.ngate.t9 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X31 iovdd.t3 sg13g2_GateDecode_0.pgate.t9 pad.t0 iovdd.t0 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X32 sg13g2_GateDecode_0.ngate.t1 a_7724_30170# iovss iovss sg13_hv_nmos ad=0.646p pd=4.48u as=0.646p ps=4.48u w=1.9u l=0.45u
X33 vdd.t6 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t2 a_8358_31526# vdd.t5 sg13_lv_pmos ad=1.615p pd=10.18u as=1.615p ps=10.18u w=4.75u l=0.13u
X34 iovss a_8358_31526# a_8358_30206# iovss sg13_hv_nmos ad=0.361p pd=2.28u as=0.646p ps=4.48u w=1.9u l=0.45u
X35 pad.t12 sg13g2_GateDecode_0.pgate.t10 iovdd.t4 iovdd.t0 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X36 pad.t1 sg13g2_GateDecode_0.pgate.t11 iovdd.t11 iovdd.t0 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X37 pad.t21 sg13g2_GateDecode_0.ngate.t10 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=2.068p ps=9.74u w=4.4u l=0.6u
X38 pad.t20 sg13g2_GateDecode_0.ngate.t11 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X39 sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq c2p_en.t1 iovss iovss sg13_lv_nmos ad=1.3362p pd=8.54u as=1.3362p ps=8.54u w=3.93u l=0.13u
X40 pad.t11 sg13g2_GateDecode_0.pgate.t12 iovdd.t2 iovdd.t0 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X41 iovdd.t16 sg13g2_GateDecode_0.pgate.t13 pad.t6 iovdd.t0 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X42 iovss sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t2 a_8358_31526# iovss sg13_lv_nmos ad=0.935p pd=6.18u as=0.935p ps=6.18u w=2.75u l=0.13u
X43 iovss sg13g2_GateDecode_0.ngate.t12 dantenna l=0.78u w=0.78u
X44 vdd.t3 c2p_en.t0 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t0 vdd.t2 sg13_lv_pmos ad=1.5876p pd=9.54u as=0.8379p ps=4.79u w=4.41u l=0.13u
X45 pad.t25 iovdd.t31 dpantenna l=1.26u w=27.78u
X46 pad.t10 sg13g2_GateDecode_0.pgate.t11 iovdd.t15 iovdd.t0 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X47 pad.t9 sg13g2_GateDecode_0.pgate.t12 iovdd.t14 iovdd.t0 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X48 iovss sg13g2_GateDecode_0.ngate.t13 pad.t19 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X49 sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq a_7750_34876# vdd.t4 sg13_lv_pmos ad=1.5876p pd=9.54u as=0.8379p ps=4.79u w=4.41u l=0.13u
X50 a_7724_30170# a_7656_30206# iovdd iovdd sg13_hv_pmos ad=0.102p pd=1.28u as=57f ps=0.68u w=0.3u l=0.45u
X51 iovdd.t13 sg13g2_GateDecode_0.pgate.t13 pad.t3 iovdd.t0 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X52 pad.t8 sg13g2_GateDecode_0.pgate.t14 iovdd.t5 iovdd.t0 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X53 iovss sg13g2_GateDecode_0.ngate.t14 pad.t17 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X54 iovss sg13g2_GateDecode_0.ngate.t15 pad.t20 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X55 sg13g2_GateDecode_0.pgate.t0 a_8426_30170# iovdd iovdd sg13_hv_pmos ad=1.326p pd=8.48u as=1.326p ps=8.48u w=3.9u l=0.45u
X56 pad.t7 sg13g2_GateDecode_0.pgate.t14 iovdd.t6 iovdd.t0 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X57 vdd.t9 sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq a_7656_31526# vdd.t5 sg13_lv_pmos ad=1.615p pd=10.18u as=1.615p ps=10.18u w=4.75u l=0.13u
X58 pad.t6 sg13g2_GateDecode_0.pgate.t15 iovdd.t12 iovdd.t0 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X59 pad.t26 iovdd.t31 dpantenna l=1.26u w=27.78u
X60 a_8230_33842# c2p.t0 iovss iovss sg13_lv_nmos ad=0.7467p pd=4.31u as=1.3362p ps=8.54u w=3.93u l=0.13u
X61 iovss a_7656_31526# a_7656_30206# iovss sg13_hv_nmos ad=0.361p pd=2.28u as=0.646p ps=4.48u w=1.9u l=0.45u
X62 iovdd.t7 sg13g2_GateDecode_0.pgate.t16 pad.t5 iovdd.t0 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X63 pad.t16 sg13g2_GateDecode_0.ngate.t16 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X64 iovss sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq a_7656_31526# iovss sg13_lv_nmos ad=0.935p pd=6.18u as=0.935p ps=6.18u w=2.75u l=0.13u
X65 a_8426_30170# sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t3 iovss iovss sg13_hv_nmos ad=0.646p pd=4.48u as=0.361p ps=2.28u w=1.9u l=0.45u
X66 iovdd a_8426_30170# a_8358_30206# iovdd sg13_hv_pmos ad=57f pd=0.68u as=0.102p ps=1.28u w=0.3u l=0.45u
X67 iovss pad.t27 dantenna l=1.26u w=27.78u
X68 sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq c2p.t1 iovss iovss sg13_lv_nmos ad=0.7467p pd=4.31u as=1.3362p ps=8.54u w=3.93u l=0.13u
X69 iovdd.t4 sg13g2_GateDecode_0.pgate.t16 pad.t4 iovdd.t0 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X70 pad.t3 sg13g2_GateDecode_0.pgate.t15 iovdd.t3 iovdd.t0 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X71 pad.t2 sg13g2_GateDecode_0.pgate.t17 iovdd.t8 iovdd.t0 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X72 sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq c2p_en.t1 vdd.t1 vdd.t0 sg13_lv_pmos ad=1.4994p pd=9.5u as=1.4994p ps=9.5u w=4.41u l=0.13u
X73 sg13g2_GateDecode_0.pgate.t1 a_8426_30170# iovss iovss sg13_hv_nmos ad=0.646p pd=4.48u as=0.646p ps=4.48u w=1.9u l=0.45u
X74 iovdd.t2 sg13g2_GateDecode_0.pgate.t3 pad.t1 iovdd.t0 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X75 pad.t22 sg13g2_GateDecode_0.ngate.t17 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X76 pad.t0 sg13g2_GateDecode_0.pgate.t17 iovdd.t1 iovdd.t0 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
R0 sg13g2_GateDecode_0.sg13g2_LevelUp_1.o sg13g2_GateDecode_0.pgate.n19 38.7086
R1 sg13g2_GateDecode_0.pgate.t0 sg13g2_GateDecode_0.pgate.n0 17.0005
R2 sg13g2_GateDecode_0.pgate.n18 sg13g2_GateDecode_0.pgate.n16 9.58949
R3 sg13g2_GateDecode_0.pgate.n17 sg13g2_GateDecode_0.pgate.n2 9.00605
R4 sg13g2_GateDecode_0.pgate.n19 sg13g2_GateDecode_0.pgate.n18 9.0005
R5 sg13g2_GateDecode_0.pgate.n3 sg13g2_GateDecode_0.pgate.t7 7.94005
R6 sg13g2_GateDecode_0.pgate.n16 sg13g2_GateDecode_0.pgate.t5 7.08755
R7 sg13g2_GateDecode_0.pgate.n3 sg13g2_GateDecode_0.pgate.t13 7.08755
R8 sg13g2_GateDecode_0.pgate.n4 sg13g2_GateDecode_0.pgate.t15 7.08755
R9 sg13g2_GateDecode_0.pgate.n5 sg13g2_GateDecode_0.pgate.t9 7.08755
R10 sg13g2_GateDecode_0.pgate.n6 sg13g2_GateDecode_0.pgate.t17 7.08755
R11 sg13g2_GateDecode_0.pgate.n7 sg13g2_GateDecode_0.pgate.t6 7.08755
R12 sg13g2_GateDecode_0.pgate.n8 sg13g2_GateDecode_0.pgate.t14 7.08755
R13 sg13g2_GateDecode_0.pgate.n9 sg13g2_GateDecode_0.pgate.t8 7.08755
R14 sg13g2_GateDecode_0.pgate.n10 sg13g2_GateDecode_0.pgate.t12 7.08755
R15 sg13g2_GateDecode_0.pgate.n11 sg13g2_GateDecode_0.pgate.t3 7.08755
R16 sg13g2_GateDecode_0.pgate.n12 sg13g2_GateDecode_0.pgate.t11 7.08755
R17 sg13g2_GateDecode_0.pgate.n13 sg13g2_GateDecode_0.pgate.t4 7.08755
R18 sg13g2_GateDecode_0.pgate.n14 sg13g2_GateDecode_0.pgate.t10 7.08755
R19 sg13g2_GateDecode_0.pgate.n15 sg13g2_GateDecode_0.pgate.t16 7.08755
R20 sg13g2_GateDecode_0.pgate.n0 sg13g2_GateDecode_0.pgate.t1 4.53355
R21 sg13g2_GateDecode_0.pgate.n17 sg13g2_GateDecode_0.pgate.t2 4.2615
R22 sg13g2_GateDecode_0.pgate.n1 sg13g2_GateDecode_0.pgate.t0 2.28308
R23 sg13g2_GateDecode_0.sg13g2_LevelUp_1.o sg13g2_GateDecode_0.pgate.n1 1.9798
R24 sg13g2_GateDecode_0.pgate.n4 sg13g2_GateDecode_0.pgate.n3 1.22425
R25 sg13g2_GateDecode_0.pgate.n6 sg13g2_GateDecode_0.pgate.n5 1.22425
R26 sg13g2_GateDecode_0.pgate.n8 sg13g2_GateDecode_0.pgate.n7 1.22425
R27 sg13g2_GateDecode_0.pgate.n10 sg13g2_GateDecode_0.pgate.n9 1.22425
R28 sg13g2_GateDecode_0.pgate.n12 sg13g2_GateDecode_0.pgate.n11 1.22425
R29 sg13g2_GateDecode_0.pgate.n14 sg13g2_GateDecode_0.pgate.n13 1.22425
R30 sg13g2_GateDecode_0.pgate.n16 sg13g2_GateDecode_0.pgate.n15 1.22425
R31 sg13g2_GateDecode_0.pgate.n5 sg13g2_GateDecode_0.pgate.n4 0.853
R32 sg13g2_GateDecode_0.pgate.n7 sg13g2_GateDecode_0.pgate.n6 0.853
R33 sg13g2_GateDecode_0.pgate.n9 sg13g2_GateDecode_0.pgate.n8 0.853
R34 sg13g2_GateDecode_0.pgate.n11 sg13g2_GateDecode_0.pgate.n10 0.853
R35 sg13g2_GateDecode_0.pgate.n13 sg13g2_GateDecode_0.pgate.n12 0.853
R36 sg13g2_GateDecode_0.pgate.n15 sg13g2_GateDecode_0.pgate.n14 0.853
R37 sg13g2_GateDecode_0.pgate.n19 sg13g2_GateDecode_0.pgate.n2 0.2117
R38 sg13g2_GateDecode_0.pgate.n18 sg13g2_GateDecode_0.pgate.n17 0.201404
R39 sg13g2_GateDecode_0.pgate.n2 sg13g2_Clamp_P15N15D_0.gate 0.0841
R40 sg13g2_GateDecode_0.pgate.n1 sg13g2_GateDecode_0.pgate.n0 0.0738333
R41 iovdd.n305 iovdd.n304 10.8089
R42 iovdd.n299 iovdd.n298 10.8089
R43 iovdd.n268 iovdd.n267 10.8089
R44 iovdd.n244 iovdd.n243 10.8089
R45 iovdd.n241 iovdd.n240 10.8089
R46 iovdd.n271 iovdd.n270 10.8089
R47 iovdd.n302 iovdd.n120 10.8089
R48 iovdd.n264 iovdd.n263 10.8089
R49 iovdd.n277 iovdd.n276 9.0005
R50 iovdd.n445 iovdd.n444 9.0005
R51 iovdd.n442 iovdd.n441 9.0005
R52 iovdd.n427 iovdd.n426 9.0005
R53 iovdd.n236 iovdd.n30 9.0005
R54 iovdd.n468 iovdd.n467 9.0005
R55 iovdd.n424 iovdd.n423 9.0005
R56 iovdd.n465 iovdd.n464 9.0005
R57 iovdd.n500 iovdd.n31 5.66717
R58 iovdd.n501 iovdd.n500 5.66717
R59 iovdd.n457 iovdd.n456 5.66717
R60 iovdd.n456 iovdd.n455 5.66717
R61 iovdd.n437 iovdd.n111 5.66717
R62 iovdd.n438 iovdd.n437 5.66717
R63 iovdd.n419 iovdd.n407 5.66717
R64 iovdd.n420 iovdd.n419 5.66717
R65 iovdd.n415 iovdd.n414 5.66717
R66 iovdd.n414 iovdd.n413 5.66717
R67 iovdd.n430 iovdd.n428 4.9805
R68 iovdd.n104 iovdd.n102 4.9805
R69 iovdd.n448 iovdd.n446 4.9805
R70 iovdd.n471 iovdd.n469 4.9805
R71 iovdd.n506 iovdd.n505 4.9805
R72 iovdd.n274 iovdd.n272 4.9805
R73 iovdd.n80 iovdd.n78 4.9805
R74 iovdd.n509 iovdd.n21 4.28068
R75 iovdd.n511 iovdd.n18 4.2505
R76 iovdd.n398 iovdd.n396 3.0005
R77 iovdd.n400 iovdd.n395 3.0005
R78 iovdd.n430 iovdd.n429 3.0005
R79 iovdd.n104 iovdd.n103 3.0005
R80 iovdd.n448 iovdd.n447 3.0005
R81 iovdd.n274 iovdd.n273 3.0005
R82 iovdd.n471 iovdd.n470 3.0005
R83 iovdd.n505 iovdd.n504 3.0005
R84 iovdd.n422 iovdd.n421 3.0005
R85 iovdd.n432 iovdd.n431 3.0005
R86 iovdd.n440 iovdd.n439 3.0005
R87 iovdd.n450 iovdd.n449 3.0005
R88 iovdd.n275 iovdd.n91 3.0005
R89 iovdd.n473 iovdd.n472 3.0005
R90 iovdd.n503 iovdd.n502 3.0005
R91 iovdd.n463 iovdd.n462 3.0005
R92 iovdd.n80 iovdd.n79 3.0005
R93 iovdd.t31 iovdd.n498 2.83433
R94 iovdd.t31 iovdd.n483 2.83433
R95 iovdd.t31 iovdd.n482 2.83433
R96 iovdd.t31 iovdd.n481 2.83433
R97 iovdd.t31 iovdd.n480 2.83433
R98 iovdd.t31 iovdd.n479 2.83433
R99 iovdd.t31 iovdd.n33 2.83433
R100 iovdd.n499 iovdd.t31 2.83433
R101 iovdd.t31 iovdd.n478 2.83433
R102 iovdd.t31 iovdd.n68 2.83433
R103 iovdd.t31 iovdd.n67 2.83433
R104 iovdd.t31 iovdd.n66 2.83433
R105 iovdd.t31 iovdd.n65 2.83433
R106 iovdd.t31 iovdd.n64 2.83433
R107 iovdd.t31 iovdd.n63 2.83433
R108 iovdd.t31 iovdd.n62 2.83433
R109 iovdd.t31 iovdd.n61 2.83433
R110 iovdd.t31 iovdd.n60 2.83433
R111 iovdd.t31 iovdd.n59 2.83433
R112 iovdd.t31 iovdd.n58 2.83433
R113 iovdd.t31 iovdd.n57 2.83433
R114 iovdd.t31 iovdd.n56 2.83433
R115 iovdd.t31 iovdd.n55 2.83433
R116 iovdd.t31 iovdd.n54 2.83433
R117 iovdd.t31 iovdd.n53 2.83433
R118 iovdd.t31 iovdd.n52 2.83433
R119 iovdd.t31 iovdd.n51 2.83433
R120 iovdd.t31 iovdd.n50 2.83433
R121 iovdd.t31 iovdd.n49 2.83433
R122 iovdd.t31 iovdd.n48 2.83433
R123 iovdd.t31 iovdd.n47 2.83433
R124 iovdd.t31 iovdd.n46 2.83433
R125 iovdd.t31 iovdd.n45 2.83433
R126 iovdd.t31 iovdd.n44 2.83433
R127 iovdd.t31 iovdd.n43 2.83433
R128 iovdd.t31 iovdd.n42 2.83433
R129 iovdd.t31 iovdd.n41 2.83433
R130 iovdd.t31 iovdd.n40 2.83433
R131 iovdd.t31 iovdd.n39 2.83433
R132 iovdd.t31 iovdd.n38 2.83433
R133 iovdd.t31 iovdd.n37 2.83433
R134 iovdd.t31 iovdd.n36 2.83433
R135 iovdd.n497 iovdd.n496 2.82693
R136 iovdd.n495 iovdd.n484 2.82693
R137 iovdd.n494 iovdd.n485 2.82693
R138 iovdd.n493 iovdd.n486 2.82693
R139 iovdd.n492 iovdd.n487 2.82693
R140 iovdd.n491 iovdd.n488 2.82693
R141 iovdd.n490 iovdd.n489 2.82693
R142 iovdd.n34 iovdd.n32 2.82693
R143 iovdd.n477 iovdd.n476 2.82693
R144 iovdd.n475 iovdd.n69 2.82693
R145 iovdd.n474 iovdd.n70 2.82693
R146 iovdd.n72 iovdd.n71 2.82693
R147 iovdd.n82 iovdd.n81 2.82693
R148 iovdd.n84 iovdd.n83 2.82693
R149 iovdd.n86 iovdd.n85 2.82693
R150 iovdd.n461 iovdd.n87 2.82693
R151 iovdd.n460 iovdd.n88 2.82693
R152 iovdd.n459 iovdd.n89 2.82693
R153 iovdd.n458 iovdd.n90 2.82693
R154 iovdd.n454 iovdd.n92 2.82693
R155 iovdd.n453 iovdd.n93 2.82693
R156 iovdd.n452 iovdd.n94 2.82693
R157 iovdd.n451 iovdd.n95 2.82693
R158 iovdd.n97 iovdd.n96 2.82693
R159 iovdd.n106 iovdd.n105 2.82693
R160 iovdd.n108 iovdd.n107 2.82693
R161 iovdd.n110 iovdd.n109 2.82693
R162 iovdd.n436 iovdd.n112 2.82693
R163 iovdd.n435 iovdd.n113 2.82693
R164 iovdd.n434 iovdd.n114 2.82693
R165 iovdd.n433 iovdd.n115 2.82693
R166 iovdd.n117 iovdd.n116 2.82693
R167 iovdd.n402 iovdd.n401 2.82693
R168 iovdd.n404 iovdd.n403 2.82693
R169 iovdd.n406 iovdd.n405 2.82693
R170 iovdd.n418 iovdd.n408 2.82693
R171 iovdd.n417 iovdd.n409 2.82693
R172 iovdd.n416 iovdd.n410 2.82693
R173 iovdd.n511 iovdd.n2 2.41731
R174 iovdd.n512 iovdd.n511 2.1192
R175 iovdd.n511 iovdd.n15 2.11861
R176 iovdd.n100 iovdd.n75 1.98828
R177 iovdd.n300 iovdd.n75 1.98792
R178 iovdd.n431 iovdd.n430 1.9805
R179 iovdd.n440 iovdd.n104 1.9805
R180 iovdd.n449 iovdd.n448 1.9805
R181 iovdd.n472 iovdd.n471 1.9805
R182 iovdd.n505 iovdd.n503 1.9805
R183 iovdd.n275 iovdd.n274 1.9805
R184 iovdd.n463 iovdd.n80 1.9805
R185 iovdd.t31 iovdd.n35 1.89
R186 iovdd.n431 iovdd.n427 1.8749
R187 iovdd.n441 iovdd.n440 1.8749
R188 iovdd.n449 iovdd.n445 1.8749
R189 iovdd.n472 iovdd.n468 1.8749
R190 iovdd.n503 iovdd.n30 1.8749
R191 iovdd.n277 iovdd.n275 1.8749
R192 iovdd.n464 iovdd.n463 1.8749
R193 iovdd.n427 iovdd.n118 1.8089
R194 iovdd.n441 iovdd.n101 1.8089
R195 iovdd.n445 iovdd.n98 1.8089
R196 iovdd.n468 iovdd.n73 1.8089
R197 iovdd.n238 iovdd.n30 1.8089
R198 iovdd.n278 iovdd.n277 1.8089
R199 iovdd.n423 iovdd.n393 1.8089
R200 iovdd.n464 iovdd.n77 1.8089
R201 iovdd.n263 iovdd.t1 1.76518
R202 iovdd.n77 iovdd.t8 1.76518
R203 iovdd.n271 iovdd.t6 1.76518
R204 iovdd.n278 iovdd.t5 1.76518
R205 iovdd.n305 iovdd.t4 1.76518
R206 iovdd.n118 iovdd.t7 1.76518
R207 iovdd.n298 iovdd.t15 1.76518
R208 iovdd.n101 iovdd.t11 1.76518
R209 iovdd.n267 iovdd.t14 1.76518
R210 iovdd.n98 iovdd.t2 1.76518
R211 iovdd.n244 iovdd.t3 1.76518
R212 iovdd.n73 iovdd.t12 1.76518
R213 iovdd.n240 iovdd.t13 1.76518
R214 iovdd.n238 iovdd.t16 1.76518
R215 iovdd.n120 iovdd.t25 1.76484
R216 iovdd.n393 iovdd.t28 1.76484
R217 iovdd.n425 iovdd.n75 1.73634
R218 iovdd.n99 iovdd.n75 1.73634
R219 iovdd.n466 iovdd.n75 1.73634
R220 iovdd.n443 iovdd.n75 1.73611
R221 iovdd.n76 iovdd.n75 1.73611
R222 iovdd.n75 iovdd.n74 1.73611
R223 iovdd.n133 iovdd.n75 1.73611
R224 iovdd.n265 iovdd.n75 1.73611
R225 iovdd.n242 iovdd.n75 1.73611
R226 iovdd.n303 iovdd.n75 1.73595
R227 iovdd.n269 iovdd.n75 1.73595
R228 iovdd.n144 iovdd.n75 1.73595
R229 iovdd.t31 iovdd.n1 1.70106
R230 iovdd.n412 iovdd.n411 1.68243
R231 iovdd.n423 iovdd.n422 1.60815
R232 iovdd.n306 iovdd.n305 1.5625
R233 iovdd.n306 iovdd.n118 1.5625
R234 iovdd.n298 iovdd.n297 1.5625
R235 iovdd.n297 iovdd.n101 1.5625
R236 iovdd.n267 iovdd.n266 1.5625
R237 iovdd.n266 iovdd.n98 1.5625
R238 iovdd.n245 iovdd.n244 1.5625
R239 iovdd.n245 iovdd.n73 1.5625
R240 iovdd.n240 iovdd.n239 1.5625
R241 iovdd.n239 iovdd.n238 1.5625
R242 iovdd.n279 iovdd.n271 1.5625
R243 iovdd.n279 iovdd.n278 1.5625
R244 iovdd.n392 iovdd.n120 1.5625
R245 iovdd.n393 iovdd.n392 1.5625
R246 iovdd.n263 iovdd.n262 1.5625
R247 iovdd.n262 iovdd.n77 1.5625
R248 iovdd iovdd.n119 1.43219
R249 iovdd.n241 iovdd.n237 1.42534
R250 iovdd.n237 iovdd.n236 1.42433
R251 iovdd.n301 iovdd 1.39634
R252 iovdd.n424 iovdd.n119 1.33976
R253 iovdd.n302 iovdd.n301 1.33311
R254 iovdd.n511 iovdd.n14 1.28534
R255 iovdd.n511 iovdd.n20 1.28534
R256 iovdd.n355 iovdd.n351 0.826084
R257 iovdd.n188 iovdd.n181 0.826084
R258 iovdd.n358 iovdd.n350 0.818682
R259 iovdd.n349 iovdd.n342 0.818682
R260 iovdd.n365 iovdd.n341 0.818682
R261 iovdd.n366 iovdd.n340 0.818682
R262 iovdd.n339 iovdd.n332 0.818682
R263 iovdd.n373 iovdd.n331 0.818682
R264 iovdd.n374 iovdd.n330 0.818682
R265 iovdd.n329 iovdd.n322 0.818682
R266 iovdd.n381 iovdd.n321 0.818682
R267 iovdd.n382 iovdd.n320 0.818682
R268 iovdd.n124 iovdd.n122 0.818682
R269 iovdd.n390 iovdd.n389 0.818682
R270 iovdd.n123 iovdd.n121 0.818682
R271 iovdd.n309 iovdd.n308 0.818682
R272 iovdd.n132 iovdd.n131 0.818682
R273 iovdd.n295 iovdd.n294 0.818682
R274 iovdd.n281 iovdd.n135 0.818682
R275 iovdd.n283 iovdd.n282 0.818682
R276 iovdd.n143 iovdd.n142 0.818682
R277 iovdd.n260 iovdd.n259 0.818682
R278 iovdd.n146 iovdd.n145 0.818682
R279 iovdd.n248 iovdd.n247 0.818682
R280 iovdd.n234 iovdd.n153 0.818682
R281 iovdd.n233 iovdd.n232 0.818682
R282 iovdd.n155 iovdd.n154 0.818682
R283 iovdd.n221 iovdd.n220 0.818682
R284 iovdd.n219 iovdd.n162 0.818682
R285 iovdd.n218 iovdd.n217 0.818682
R286 iovdd.n164 iovdd.n163 0.818682
R287 iovdd.n206 iovdd.n205 0.818682
R288 iovdd.n204 iovdd.n171 0.818682
R289 iovdd.n203 iovdd.n202 0.818682
R290 iovdd.n173 iovdd.n172 0.818682
R291 iovdd.n191 iovdd.n190 0.818682
R292 iovdd.n189 iovdd.n180 0.818682
R293 iovdd.n187 iovdd.n186 0.818682
R294 iovdd.n182 iovdd.n180 0.818682
R295 iovdd.n192 iovdd.n191 0.818682
R296 iovdd.n193 iovdd.n173 0.818682
R297 iovdd.n202 iovdd.n201 0.818682
R298 iovdd.n175 iovdd.n171 0.818682
R299 iovdd.n207 iovdd.n206 0.818682
R300 iovdd.n208 iovdd.n164 0.818682
R301 iovdd.n217 iovdd.n216 0.818682
R302 iovdd.n166 iovdd.n162 0.818682
R303 iovdd.n222 iovdd.n221 0.818682
R304 iovdd.n223 iovdd.n155 0.818682
R305 iovdd.n232 iovdd.n231 0.818682
R306 iovdd.n157 iovdd.n153 0.818682
R307 iovdd.n249 iovdd.n248 0.818682
R308 iovdd.n250 iovdd.n146 0.818682
R309 iovdd.n259 iovdd.n258 0.818682
R310 iovdd.n148 iovdd.n142 0.818682
R311 iovdd.n284 iovdd.n283 0.818682
R312 iovdd.n285 iovdd.n135 0.818682
R313 iovdd.n294 iovdd.n293 0.818682
R314 iovdd.n137 iovdd.n131 0.818682
R315 iovdd.n310 iovdd.n309 0.818682
R316 iovdd.n311 iovdd.n123 0.818682
R317 iovdd.n389 iovdd.n388 0.818682
R318 iovdd.n126 iovdd.n124 0.818682
R319 iovdd.n383 iovdd.n382 0.818682
R320 iovdd.n381 iovdd.n380 0.818682
R321 iovdd.n323 iovdd.n322 0.818682
R322 iovdd.n375 iovdd.n374 0.818682
R323 iovdd.n373 iovdd.n372 0.818682
R324 iovdd.n333 iovdd.n332 0.818682
R325 iovdd.n367 iovdd.n366 0.818682
R326 iovdd.n365 iovdd.n364 0.818682
R327 iovdd.n343 iovdd.n342 0.818682
R328 iovdd.n359 iovdd.n358 0.818682
R329 iovdd.n357 iovdd.n356 0.818682
R330 iovdd.n511 iovdd.n22 0.671789
R331 iovdd.n511 iovdd.n6 0.671602
R332 iovdd.n511 iovdd.n28 0.671602
R333 iovdd.n511 iovdd.n12 0.671423
R334 iovdd.n511 iovdd.n24 0.588672
R335 iovdd.n511 iovdd.n26 0.588672
R336 iovdd.n511 iovdd.n29 0.588672
R337 iovdd.n511 iovdd.n11 0.588437
R338 iovdd.n511 iovdd.n9 0.588437
R339 iovdd.n511 iovdd.n7 0.588437
R340 iovdd.n511 iovdd.n23 0.588437
R341 iovdd.n511 iovdd.n25 0.588437
R342 iovdd.n511 iovdd.n27 0.588437
R343 iovdd.n511 iovdd.n10 0.588281
R344 iovdd.n511 iovdd.n8 0.588281
R345 iovdd.n511 iovdd.n5 0.588281
R346 iovdd.n511 iovdd.n3 0.588266
R347 iovdd.n444 iovdd.n443 0.515695
R348 iovdd.n268 iovdd.n133 0.515695
R349 iovdd.n425 iovdd.n424 0.513735
R350 iovdd.n303 iovdd.n302 0.513312
R351 iovdd.n511 iovdd.n510 0.503491
R352 iovdd.n270 iovdd.n269 0.502871
R353 iovdd.n276 iovdd.n99 0.502476
R354 iovdd.n511 iovdd.n17 0.502128
R355 iovdd.n465 iovdd.n76 0.489812
R356 iovdd.n265 iovdd.n264 0.489812
R357 iovdd.n467 iovdd.n74 0.481088
R358 iovdd.n243 iovdd.n242 0.481088
R359 iovdd.n300 iovdd.n299 0.479418
R360 iovdd.n442 iovdd.n100 0.479034
R361 iovdd.n426 iovdd.n100 0.477001
R362 iovdd.n243 iovdd.n144 0.476989
R363 iovdd.n304 iovdd.n300 0.476595
R364 iovdd.n467 iovdd.n466 0.476594
R365 iovdd.n466 iovdd.n465 0.468441
R366 iovdd.n264 iovdd.n144 0.468018
R367 iovdd.n236 iovdd.n74 0.46393
R368 iovdd.n242 iovdd.n241 0.46393
R369 iovdd.n276 iovdd.n76 0.455206
R370 iovdd.n270 iovdd.n265 0.455206
R371 iovdd.n444 iovdd.n99 0.442559
R372 iovdd.n269 iovdd.n268 0.442135
R373 iovdd.n304 iovdd.n303 0.431695
R374 iovdd.n426 iovdd.n425 0.4313
R375 iovdd.n443 iovdd.n442 0.429323
R376 iovdd.n299 iovdd.n133 0.429323
R377 iovdd.n189 iovdd.n188 0.416993
R378 iovdd.n351 iovdd.n350 0.416993
R379 iovdd.n507 iovdd.n506 0.328683
R380 iovdd.n508 iovdd.n507 0.270343
R381 iovdd.n508 iovdd.n4 0.258522
R382 iovdd.n511 iovdd.n4 0.254672
R383 iovdd.n398 iovdd.n397 0.2505
R384 iovdd.n400 iovdd.n399 0.2505
R385 iovdd.n422 iovdd.n394 0.2505
R386 iovdd.n504 iovdd.n4 0.227256
R387 iovdd.n183 iovdd.n181 0.201704
R388 iovdd.n355 iovdd.n354 0.2005
R389 iovdd.n348 iovdd.n347 0.2005
R390 iovdd.n361 iovdd.n360 0.2005
R391 iovdd.n363 iovdd.n362 0.2005
R392 iovdd.n338 iovdd.n337 0.2005
R393 iovdd.n369 iovdd.n368 0.2005
R394 iovdd.n371 iovdd.n370 0.2005
R395 iovdd.n328 iovdd.n327 0.2005
R396 iovdd.n377 iovdd.n376 0.2005
R397 iovdd.n379 iovdd.n378 0.2005
R398 iovdd.n319 iovdd.n318 0.2005
R399 iovdd.n385 iovdd.n384 0.2005
R400 iovdd.n387 iovdd.n386 0.2005
R401 iovdd.n127 iovdd.n125 0.2005
R402 iovdd.n313 iovdd.n312 0.2005
R403 iovdd.n130 iovdd.n129 0.2005
R404 iovdd.n292 iovdd.n291 0.2005
R405 iovdd.n138 iovdd.n136 0.2005
R406 iovdd.n287 iovdd.n286 0.2005
R407 iovdd.n141 iovdd.n140 0.2005
R408 iovdd.n257 iovdd.n256 0.2005
R409 iovdd.n149 iovdd.n147 0.2005
R410 iovdd.n252 iovdd.n251 0.2005
R411 iovdd.n152 iovdd.n151 0.2005
R412 iovdd.n230 iovdd.n229 0.2005
R413 iovdd.n158 iovdd.n156 0.2005
R414 iovdd.n225 iovdd.n224 0.2005
R415 iovdd.n161 iovdd.n160 0.2005
R416 iovdd.n215 iovdd.n214 0.2005
R417 iovdd.n167 iovdd.n165 0.2005
R418 iovdd.n210 iovdd.n209 0.2005
R419 iovdd.n170 iovdd.n169 0.2005
R420 iovdd.n200 iovdd.n199 0.2005
R421 iovdd.n176 iovdd.n174 0.2005
R422 iovdd.n195 iovdd.n194 0.2005
R423 iovdd.n179 iovdd.n178 0.2005
R424 iovdd.n185 iovdd.n184 0.2005
R425 iovdd.n262 iovdd.n261 0.191989
R426 iovdd.n280 iovdd.n279 0.191989
R427 iovdd.n266 iovdd.n134 0.191989
R428 iovdd.n297 iovdd.n296 0.191989
R429 iovdd.n307 iovdd.n306 0.191989
R430 iovdd.n392 iovdd.n391 0.191989
R431 iovdd.n239 iovdd.n235 0.191989
R432 iovdd.n246 iovdd.n245 0.191989
R433 iovdd.n17 iovdd.n16 0.156542
R434 iovdd.n510 iovdd.n508 0.153056
R435 iovdd.n3 iovdd.n0 0.144604
R436 iovdd.n504 iovdd.n5 0.143944
R437 iovdd.n506 iovdd.n29 0.14355
R438 iovdd.n272 iovdd.n27 0.142174
R439 iovdd.n273 iovdd.n7 0.142174
R440 iovdd.n16 iovdd.n3 0.139796
R441 iovdd.n446 iovdd.n26 0.138974
R442 iovdd.n447 iovdd.n8 0.138556
R443 iovdd.n102 iovdd.n25 0.13519
R444 iovdd.n103 iovdd.n9 0.13519
R445 iovdd.n429 iovdd.n11 0.135097
R446 iovdd.n428 iovdd.n23 0.135097
R447 iovdd.n470 iovdd.n6 0.133441
R448 iovdd.n469 iovdd.n28 0.133441
R449 iovdd.n428 iovdd.n24 0.13199
R450 iovdd.n103 iovdd.n10 0.131722
R451 iovdd.n78 iovdd.n28 0.131626
R452 iovdd.n79 iovdd.n6 0.131626
R453 iovdd.n429 iovdd.n10 0.131572
R454 iovdd.n102 iovdd.n24 0.131328
R455 iovdd.n396 iovdd.n23 0.128206
R456 iovdd.n395 iovdd.n11 0.128206
R457 iovdd.n447 iovdd.n9 0.128113
R458 iovdd.n446 iovdd.n25 0.128113
R459 iovdd.n510 iovdd.n509 0.127471
R460 iovdd.n395 iovdd.n12 0.124896
R461 iovdd.n273 iovdd.n8 0.124738
R462 iovdd.n19 iovdd.n17 0.124655
R463 iovdd.n396 iovdd.n22 0.124514
R464 iovdd.n272 iovdd.n26 0.124344
R465 iovdd.n79 iovdd.n7 0.121129
R466 iovdd.n78 iovdd.n27 0.121129
R467 iovdd.n469 iovdd.n29 0.119767
R468 iovdd.n470 iovdd.n5 0.11935
R469 iovdd.n397 iovdd.n22 0.117846
R470 iovdd.n399 iovdd.n12 0.117444
R471 iovdd.n354 iovdd.n353 0.1105
R472 iovdd.n352 iovdd.n347 0.1105
R473 iovdd.n361 iovdd.n346 0.1105
R474 iovdd.n362 iovdd.n345 0.1105
R475 iovdd.n344 iovdd.n337 0.1105
R476 iovdd.n369 iovdd.n336 0.1105
R477 iovdd.n370 iovdd.n335 0.1105
R478 iovdd.n334 iovdd.n327 0.1105
R479 iovdd.n377 iovdd.n326 0.1105
R480 iovdd.n378 iovdd.n325 0.1105
R481 iovdd.n324 iovdd.n318 0.1105
R482 iovdd.n385 iovdd.n317 0.1105
R483 iovdd.n386 iovdd.n316 0.1105
R484 iovdd.n315 iovdd.n127 0.1105
R485 iovdd.n314 iovdd.n313 0.1105
R486 iovdd.n129 iovdd.n128 0.1105
R487 iovdd.n291 iovdd.n290 0.1105
R488 iovdd.n289 iovdd.n138 0.1105
R489 iovdd.n288 iovdd.n287 0.1105
R490 iovdd.n140 iovdd.n139 0.1105
R491 iovdd.n256 iovdd.n255 0.1105
R492 iovdd.n254 iovdd.n149 0.1105
R493 iovdd.n253 iovdd.n252 0.1105
R494 iovdd.n151 iovdd.n150 0.1105
R495 iovdd.n229 iovdd.n228 0.1105
R496 iovdd.n227 iovdd.n158 0.1105
R497 iovdd.n226 iovdd.n225 0.1105
R498 iovdd.n160 iovdd.n159 0.1105
R499 iovdd.n214 iovdd.n213 0.1105
R500 iovdd.n212 iovdd.n167 0.1105
R501 iovdd.n211 iovdd.n210 0.1105
R502 iovdd.n169 iovdd.n168 0.1105
R503 iovdd.n199 iovdd.n198 0.1105
R504 iovdd.n197 iovdd.n176 0.1105
R505 iovdd.n196 iovdd.n195 0.1105
R506 iovdd.n178 iovdd.n177 0.1105
R507 iovdd.n511 iovdd.n507 0.0888927
R508 iovdd.n16 iovdd.n14 0.0878254
R509 iovdd.n20 iovdd.n19 0.0878254
R510 iovdd.n496 iovdd.n2 0.0776874
R511 iovdd.n422 iovdd.n400 0.0751466
R512 iovdd.n400 iovdd.n398 0.0751466
R513 iovdd.n397 iovdd.n20 0.0732046
R514 iovdd.n399 iovdd.n14 0.0732046
R515 iovdd.n413 iovdd.n412 0.0727627
R516 iovdd.n412 iovdd.n0 0.0709471
R517 iovdd.n496 iovdd.n495 0.0607875
R518 iovdd.n495 iovdd.n494 0.0607875
R519 iovdd.n494 iovdd.n493 0.0607875
R520 iovdd.n493 iovdd.n492 0.0607875
R521 iovdd.n492 iovdd.n491 0.0607875
R522 iovdd.n491 iovdd.n490 0.0607875
R523 iovdd.n476 iovdd.n32 0.0607875
R524 iovdd.n476 iovdd.n475 0.0607875
R525 iovdd.n475 iovdd.n474 0.0607875
R526 iovdd.n82 iovdd.n72 0.0607875
R527 iovdd.n84 iovdd.n82 0.0607875
R528 iovdd.n86 iovdd.n84 0.0607875
R529 iovdd.n461 iovdd.n460 0.0607875
R530 iovdd.n460 iovdd.n459 0.0607875
R531 iovdd.n459 iovdd.n458 0.0607875
R532 iovdd.n454 iovdd.n453 0.0607875
R533 iovdd.n453 iovdd.n452 0.0607875
R534 iovdd.n452 iovdd.n451 0.0607875
R535 iovdd.n106 iovdd.n97 0.0607875
R536 iovdd.n108 iovdd.n106 0.0607875
R537 iovdd.n110 iovdd.n108 0.0607875
R538 iovdd.n436 iovdd.n435 0.0607875
R539 iovdd.n435 iovdd.n434 0.0607875
R540 iovdd.n434 iovdd.n433 0.0607875
R541 iovdd.n402 iovdd.n117 0.0607875
R542 iovdd.n404 iovdd.n402 0.0607875
R543 iovdd.n406 iovdd.n404 0.0607875
R544 iovdd.n418 iovdd.n417 0.0607875
R545 iovdd.n417 iovdd.n416 0.0607875
R546 iovdd.n183 iovdd.n177 0.0568704
R547 iovdd.n509 iovdd.n2 0.0540779
R548 iovdd.t31 iovdd.n21 0.0491586
R549 iovdd.t31 iovdd.n13 0.048619
R550 iovdd.n490 iovdd.n31 0.045485
R551 iovdd.n501 iovdd.n32 0.045485
R552 iovdd.n458 iovdd.n457 0.045485
R553 iovdd.n455 iovdd.n454 0.045485
R554 iovdd.n111 iovdd.n110 0.045485
R555 iovdd.n438 iovdd.n436 0.045485
R556 iovdd.n407 iovdd.n406 0.045485
R557 iovdd.n420 iovdd.n418 0.045485
R558 iovdd.n416 iovdd.n415 0.045485
R559 iovdd.n473 iovdd.n72 0.0450485
R560 iovdd iovdd.n512 0.0429819
R561 iovdd.n462 iovdd.n86 0.0424295
R562 iovdd.n15 iovdd 0.0411071
R563 iovdd.n451 iovdd.n450 0.0354454
R564 iovdd.n432 iovdd.n117 0.0328263
R565 iovdd.n75 iovdd.t0 0.0323352
R566 iovdd.n19 iovdd.n18 0.0301825
R567 iovdd.n433 iovdd.n432 0.0284612
R568 iovdd.n502 iovdd.n501 0.026254
R569 iovdd.n450 iovdd.n97 0.0258422
R570 iovdd.n18 iovdd 0.0258175
R571 iovdd.n457 iovdd.n91 0.0236349
R572 iovdd.n421 iovdd.n420 0.0210159
R573 iovdd.n462 iovdd.n461 0.0188581
R574 iovdd.n413 iovdd.n394 0.0175238
R575 iovdd.n512 iovdd.n0 0.0169094
R576 iovdd.n439 iovdd.n111 0.0166508
R577 iovdd.n474 iovdd.n473 0.016239
R578 iovdd.n16 iovdd.n15 0.0157896
R579 iovdd.n439 iovdd.n438 0.0140317
R580 iovdd.n415 iovdd.n394 0.0131587
R581 iovdd.n421 iovdd.n407 0.00966667
R582 iovdd.n301 iovdd.n75 0.00930884
R583 iovdd.n190 iovdd.n189 0.00740196
R584 iovdd.n190 iovdd.n172 0.00740196
R585 iovdd.n203 iovdd.n172 0.00740196
R586 iovdd.n204 iovdd.n203 0.00740196
R587 iovdd.n205 iovdd.n204 0.00740196
R588 iovdd.n205 iovdd.n163 0.00740196
R589 iovdd.n218 iovdd.n163 0.00740196
R590 iovdd.n219 iovdd.n218 0.00740196
R591 iovdd.n220 iovdd.n219 0.00740196
R592 iovdd.n220 iovdd.n154 0.00740196
R593 iovdd.n233 iovdd.n154 0.00740196
R594 iovdd.n234 iovdd.n233 0.00740196
R595 iovdd.n260 iovdd.n145 0.00740196
R596 iovdd.n282 iovdd.n281 0.00740196
R597 iovdd.n308 iovdd.n132 0.00740196
R598 iovdd.n390 iovdd.n122 0.00740196
R599 iovdd.n320 iovdd.n122 0.00740196
R600 iovdd.n321 iovdd.n320 0.00740196
R601 iovdd.n329 iovdd.n321 0.00740196
R602 iovdd.n330 iovdd.n329 0.00740196
R603 iovdd.n331 iovdd.n330 0.00740196
R604 iovdd.n339 iovdd.n331 0.00740196
R605 iovdd.n340 iovdd.n339 0.00740196
R606 iovdd.n341 iovdd.n340 0.00740196
R607 iovdd.n349 iovdd.n341 0.00740196
R608 iovdd.n350 iovdd.n349 0.00740196
R609 iovdd.n187 iovdd.n180 0.00740196
R610 iovdd.n191 iovdd.n180 0.00740196
R611 iovdd.n191 iovdd.n173 0.00740196
R612 iovdd.n202 iovdd.n173 0.00740196
R613 iovdd.n202 iovdd.n171 0.00740196
R614 iovdd.n206 iovdd.n171 0.00740196
R615 iovdd.n206 iovdd.n164 0.00740196
R616 iovdd.n217 iovdd.n164 0.00740196
R617 iovdd.n217 iovdd.n162 0.00740196
R618 iovdd.n221 iovdd.n162 0.00740196
R619 iovdd.n221 iovdd.n155 0.00740196
R620 iovdd.n232 iovdd.n155 0.00740196
R621 iovdd.n232 iovdd.n153 0.00740196
R622 iovdd.n248 iovdd.n153 0.00740196
R623 iovdd.n248 iovdd.n146 0.00740196
R624 iovdd.n259 iovdd.n146 0.00740196
R625 iovdd.n259 iovdd.n142 0.00740196
R626 iovdd.n283 iovdd.n142 0.00740196
R627 iovdd.n283 iovdd.n135 0.00740196
R628 iovdd.n294 iovdd.n135 0.00740196
R629 iovdd.n294 iovdd.n131 0.00740196
R630 iovdd.n309 iovdd.n131 0.00740196
R631 iovdd.n309 iovdd.n123 0.00740196
R632 iovdd.n389 iovdd.n123 0.00740196
R633 iovdd.n389 iovdd.n124 0.00740196
R634 iovdd.n382 iovdd.n124 0.00740196
R635 iovdd.n382 iovdd.n381 0.00740196
R636 iovdd.n381 iovdd.n322 0.00740196
R637 iovdd.n374 iovdd.n322 0.00740196
R638 iovdd.n374 iovdd.n373 0.00740196
R639 iovdd.n373 iovdd.n332 0.00740196
R640 iovdd.n366 iovdd.n332 0.00740196
R641 iovdd.n366 iovdd.n365 0.00740196
R642 iovdd.n365 iovdd.n342 0.00740196
R643 iovdd.n358 iovdd.n342 0.00740196
R644 iovdd.n358 iovdd.n357 0.00740196
R645 iovdd.n455 iovdd.n91 0.00704762
R646 iovdd.n247 iovdd.n235 0.00676353
R647 iovdd.n261 iovdd.n143 0.00662549
R648 iovdd.n295 iovdd.n134 0.00648745
R649 iovdd.n307 iovdd.n121 0.00634941
R650 iovdd.n391 iovdd.n121 0.00507255
R651 iovdd.n296 iovdd.n295 0.00493451
R652 iovdd.n280 iovdd.n143 0.00479647
R653 iovdd.n247 iovdd.n246 0.00465843
R654 iovdd.n502 iovdd.n31 0.00442857
R655 iovdd.n357 iovdd.n351 0.00442211
R656 iovdd.n188 iovdd.n187 0.00442211
R657 iovdd.n119 iovdd.n75 0.00437583
R658 iovdd.n186 iovdd.n181 0.00395098
R659 iovdd.n186 iovdd.n185 0.00395098
R660 iovdd.n185 iovdd.n182 0.00395098
R661 iovdd.n182 iovdd.n179 0.00395098
R662 iovdd.n192 iovdd.n179 0.00395098
R663 iovdd.n194 iovdd.n192 0.00395098
R664 iovdd.n194 iovdd.n193 0.00395098
R665 iovdd.n193 iovdd.n174 0.00395098
R666 iovdd.n201 iovdd.n174 0.00395098
R667 iovdd.n201 iovdd.n200 0.00395098
R668 iovdd.n200 iovdd.n175 0.00395098
R669 iovdd.n175 iovdd.n170 0.00395098
R670 iovdd.n207 iovdd.n170 0.00395098
R671 iovdd.n209 iovdd.n207 0.00395098
R672 iovdd.n209 iovdd.n208 0.00395098
R673 iovdd.n208 iovdd.n165 0.00395098
R674 iovdd.n216 iovdd.n165 0.00395098
R675 iovdd.n216 iovdd.n215 0.00395098
R676 iovdd.n215 iovdd.n166 0.00395098
R677 iovdd.n166 iovdd.n161 0.00395098
R678 iovdd.n222 iovdd.n161 0.00395098
R679 iovdd.n224 iovdd.n222 0.00395098
R680 iovdd.n224 iovdd.n223 0.00395098
R681 iovdd.n223 iovdd.n156 0.00395098
R682 iovdd.n231 iovdd.n156 0.00395098
R683 iovdd.n231 iovdd.n230 0.00395098
R684 iovdd.n230 iovdd.n157 0.00395098
R685 iovdd.n157 iovdd.n152 0.00395098
R686 iovdd.n249 iovdd.n152 0.00395098
R687 iovdd.n251 iovdd.n249 0.00395098
R688 iovdd.n251 iovdd.n250 0.00395098
R689 iovdd.n250 iovdd.n147 0.00395098
R690 iovdd.n258 iovdd.n147 0.00395098
R691 iovdd.n258 iovdd.n257 0.00395098
R692 iovdd.n257 iovdd.n148 0.00395098
R693 iovdd.n148 iovdd.n141 0.00395098
R694 iovdd.n284 iovdd.n141 0.00395098
R695 iovdd.n286 iovdd.n284 0.00395098
R696 iovdd.n286 iovdd.n285 0.00395098
R697 iovdd.n285 iovdd.n136 0.00395098
R698 iovdd.n293 iovdd.n136 0.00395098
R699 iovdd.n293 iovdd.n292 0.00395098
R700 iovdd.n292 iovdd.n137 0.00395098
R701 iovdd.n137 iovdd.n130 0.00395098
R702 iovdd.n310 iovdd.n130 0.00395098
R703 iovdd.n312 iovdd.n310 0.00395098
R704 iovdd.n312 iovdd.n311 0.00395098
R705 iovdd.n311 iovdd.n125 0.00395098
R706 iovdd.n388 iovdd.n125 0.00395098
R707 iovdd.n388 iovdd.n387 0.00395098
R708 iovdd.n387 iovdd.n126 0.00395098
R709 iovdd.n384 iovdd.n126 0.00395098
R710 iovdd.n384 iovdd.n383 0.00395098
R711 iovdd.n383 iovdd.n319 0.00395098
R712 iovdd.n380 iovdd.n319 0.00395098
R713 iovdd.n380 iovdd.n379 0.00395098
R714 iovdd.n379 iovdd.n323 0.00395098
R715 iovdd.n376 iovdd.n323 0.00395098
R716 iovdd.n376 iovdd.n375 0.00395098
R717 iovdd.n375 iovdd.n328 0.00395098
R718 iovdd.n372 iovdd.n328 0.00395098
R719 iovdd.n372 iovdd.n371 0.00395098
R720 iovdd.n371 iovdd.n333 0.00395098
R721 iovdd.n368 iovdd.n333 0.00395098
R722 iovdd.n368 iovdd.n367 0.00395098
R723 iovdd.n367 iovdd.n338 0.00395098
R724 iovdd.n364 iovdd.n338 0.00395098
R725 iovdd.n364 iovdd.n363 0.00395098
R726 iovdd.n363 iovdd.n343 0.00395098
R727 iovdd.n360 iovdd.n343 0.00395098
R728 iovdd.n360 iovdd.n359 0.00395098
R729 iovdd.n359 iovdd.n348 0.00395098
R730 iovdd.n356 iovdd.n348 0.00395098
R731 iovdd.n356 iovdd.n355 0.00395098
R732 iovdd.n246 iovdd.n145 0.00324353
R733 iovdd.n282 iovdd.n280 0.00310549
R734 iovdd.n296 iovdd.n132 0.00296745
R735 iovdd.n391 iovdd.n390 0.00282941
R736 iovdd.n354 iovdd 0.00261765
R737 iovdd.n353 iovdd 0.00196667
R738 iovdd.n184 iovdd.n178 0.00191176
R739 iovdd.n195 iovdd.n178 0.00191176
R740 iovdd.n195 iovdd.n176 0.00191176
R741 iovdd.n199 iovdd.n176 0.00191176
R742 iovdd.n199 iovdd.n169 0.00191176
R743 iovdd.n210 iovdd.n169 0.00191176
R744 iovdd.n210 iovdd.n167 0.00191176
R745 iovdd.n214 iovdd.n167 0.00191176
R746 iovdd.n214 iovdd.n160 0.00191176
R747 iovdd.n225 iovdd.n160 0.00191176
R748 iovdd.n225 iovdd.n158 0.00191176
R749 iovdd.n229 iovdd.n158 0.00191176
R750 iovdd.n229 iovdd.n151 0.00191176
R751 iovdd.n252 iovdd.n151 0.00191176
R752 iovdd.n252 iovdd.n149 0.00191176
R753 iovdd.n256 iovdd.n149 0.00191176
R754 iovdd.n256 iovdd.n140 0.00191176
R755 iovdd.n287 iovdd.n140 0.00191176
R756 iovdd.n287 iovdd.n138 0.00191176
R757 iovdd.n291 iovdd.n138 0.00191176
R758 iovdd.n291 iovdd.n129 0.00191176
R759 iovdd.n313 iovdd.n129 0.00191176
R760 iovdd.n313 iovdd.n127 0.00191176
R761 iovdd.n386 iovdd.n127 0.00191176
R762 iovdd.n386 iovdd.n385 0.00191176
R763 iovdd.n385 iovdd.n318 0.00191176
R764 iovdd.n378 iovdd.n318 0.00191176
R765 iovdd.n378 iovdd.n377 0.00191176
R766 iovdd.n377 iovdd.n327 0.00191176
R767 iovdd.n370 iovdd.n327 0.00191176
R768 iovdd.n370 iovdd.n369 0.00191176
R769 iovdd.n369 iovdd.n337 0.00191176
R770 iovdd.n362 iovdd.n337 0.00191176
R771 iovdd.n362 iovdd.n361 0.00191176
R772 iovdd.n361 iovdd.n347 0.00191176
R773 iovdd.n354 iovdd.n347 0.00191176
R774 iovdd.n497 iovdd.n1 0.00170001
R775 iovdd.n184 iovdd.n183 0.0016983
R776 iovdd.n414 iovdd.n35 0.00166668
R777 iovdd.n308 iovdd.n307 0.00155255
R778 iovdd.n196 iovdd.n177 0.00147778
R779 iovdd.n197 iovdd.n196 0.00147778
R780 iovdd.n198 iovdd.n197 0.00147778
R781 iovdd.n198 iovdd.n168 0.00147778
R782 iovdd.n211 iovdd.n168 0.00147778
R783 iovdd.n212 iovdd.n211 0.00147778
R784 iovdd.n213 iovdd.n212 0.00147778
R785 iovdd.n213 iovdd.n159 0.00147778
R786 iovdd.n226 iovdd.n159 0.00147778
R787 iovdd.n227 iovdd.n226 0.00147778
R788 iovdd.n228 iovdd.n227 0.00147778
R789 iovdd.n228 iovdd.n150 0.00147778
R790 iovdd.n253 iovdd.n150 0.00147778
R791 iovdd.n254 iovdd.n253 0.00147778
R792 iovdd.n255 iovdd.n254 0.00147778
R793 iovdd.n255 iovdd.n139 0.00147778
R794 iovdd.n288 iovdd.n139 0.00147778
R795 iovdd.n289 iovdd.n288 0.00147778
R796 iovdd.n290 iovdd.n289 0.00147778
R797 iovdd.n290 iovdd.n128 0.00147778
R798 iovdd.n314 iovdd.n128 0.00147778
R799 iovdd.n315 iovdd.n314 0.00147778
R800 iovdd.n316 iovdd.n315 0.00147778
R801 iovdd.n317 iovdd.n316 0.00147778
R802 iovdd.n324 iovdd.n317 0.00147778
R803 iovdd.n325 iovdd.n324 0.00147778
R804 iovdd.n326 iovdd.n325 0.00147778
R805 iovdd.n334 iovdd.n326 0.00147778
R806 iovdd.n335 iovdd.n334 0.00147778
R807 iovdd.n336 iovdd.n335 0.00147778
R808 iovdd.n344 iovdd.n336 0.00147778
R809 iovdd.n345 iovdd.n344 0.00147778
R810 iovdd.n346 iovdd.n345 0.00147778
R811 iovdd.n352 iovdd.n346 0.00147778
R812 iovdd.n353 iovdd.n352 0.00147778
R813 iovdd.n281 iovdd.n134 0.00141451
R814 iovdd.n411 iovdd.n35 0.00133329
R815 iovdd.n511 iovdd.n1 0.00129996
R816 iovdd.n261 iovdd.n260 0.00127647
R817 iovdd.n235 iovdd.n234 0.00113843
R818 iovdd.n237 iovdd.n75 0.00100275
R819 iovdd.n511 iovdd.n13 0.001
R820 iovdd.n511 iovdd.n21 0.001
R821 iovdd.n498 iovdd.n484 0.001
R822 iovdd.n485 iovdd.n483 0.001
R823 iovdd.n486 iovdd.n482 0.001
R824 iovdd.n487 iovdd.n481 0.001
R825 iovdd.n488 iovdd.n480 0.001
R826 iovdd.n489 iovdd.n479 0.001
R827 iovdd.n500 iovdd.n33 0.001
R828 iovdd.n499 iovdd.n34 0.001
R829 iovdd.n478 iovdd.n477 0.001
R830 iovdd.n69 iovdd.n68 0.001
R831 iovdd.n70 iovdd.n67 0.001
R832 iovdd.n71 iovdd.n66 0.001
R833 iovdd.n81 iovdd.n65 0.001
R834 iovdd.n83 iovdd.n64 0.001
R835 iovdd.n85 iovdd.n63 0.001
R836 iovdd.n87 iovdd.n62 0.001
R837 iovdd.n88 iovdd.n61 0.001
R838 iovdd.n89 iovdd.n60 0.001
R839 iovdd.n90 iovdd.n59 0.001
R840 iovdd.n456 iovdd.n58 0.001
R841 iovdd.n92 iovdd.n57 0.001
R842 iovdd.n93 iovdd.n56 0.001
R843 iovdd.n94 iovdd.n55 0.001
R844 iovdd.n95 iovdd.n54 0.001
R845 iovdd.n96 iovdd.n53 0.001
R846 iovdd.n105 iovdd.n52 0.001
R847 iovdd.n107 iovdd.n51 0.001
R848 iovdd.n109 iovdd.n50 0.001
R849 iovdd.n437 iovdd.n49 0.001
R850 iovdd.n112 iovdd.n48 0.001
R851 iovdd.n113 iovdd.n47 0.001
R852 iovdd.n114 iovdd.n46 0.001
R853 iovdd.n115 iovdd.n45 0.001
R854 iovdd.n116 iovdd.n44 0.001
R855 iovdd.n401 iovdd.n43 0.001
R856 iovdd.n403 iovdd.n42 0.001
R857 iovdd.n405 iovdd.n41 0.001
R858 iovdd.n419 iovdd.n40 0.001
R859 iovdd.n408 iovdd.n39 0.001
R860 iovdd.n409 iovdd.n38 0.001
R861 iovdd.n410 iovdd.n37 0.001
R862 iovdd.n414 iovdd.n36 0.001
R863 iovdd.n411 iovdd.n13 0.001
R864 iovdd.n498 iovdd.n497 0.001
R865 iovdd.n484 iovdd.n483 0.001
R866 iovdd.n485 iovdd.n482 0.001
R867 iovdd.n486 iovdd.n481 0.001
R868 iovdd.n487 iovdd.n480 0.001
R869 iovdd.n488 iovdd.n479 0.001
R870 iovdd.n489 iovdd.n33 0.001
R871 iovdd.n500 iovdd.n499 0.001
R872 iovdd.n478 iovdd.n34 0.001
R873 iovdd.n477 iovdd.n68 0.001
R874 iovdd.n69 iovdd.n67 0.001
R875 iovdd.n70 iovdd.n66 0.001
R876 iovdd.n71 iovdd.n65 0.001
R877 iovdd.n81 iovdd.n64 0.001
R878 iovdd.n83 iovdd.n63 0.001
R879 iovdd.n85 iovdd.n62 0.001
R880 iovdd.n87 iovdd.n61 0.001
R881 iovdd.n88 iovdd.n60 0.001
R882 iovdd.n89 iovdd.n59 0.001
R883 iovdd.n90 iovdd.n58 0.001
R884 iovdd.n456 iovdd.n57 0.001
R885 iovdd.n92 iovdd.n56 0.001
R886 iovdd.n93 iovdd.n55 0.001
R887 iovdd.n94 iovdd.n54 0.001
R888 iovdd.n95 iovdd.n53 0.001
R889 iovdd.n96 iovdd.n52 0.001
R890 iovdd.n105 iovdd.n51 0.001
R891 iovdd.n107 iovdd.n50 0.001
R892 iovdd.n109 iovdd.n49 0.001
R893 iovdd.n437 iovdd.n48 0.001
R894 iovdd.n112 iovdd.n47 0.001
R895 iovdd.n113 iovdd.n46 0.001
R896 iovdd.n114 iovdd.n45 0.001
R897 iovdd.n115 iovdd.n44 0.001
R898 iovdd.n116 iovdd.n43 0.001
R899 iovdd.n401 iovdd.n42 0.001
R900 iovdd.n403 iovdd.n41 0.001
R901 iovdd.n405 iovdd.n40 0.001
R902 iovdd.n419 iovdd.n39 0.001
R903 iovdd.n408 iovdd.n38 0.001
R904 iovdd.n409 iovdd.n37 0.001
R905 iovdd.n410 iovdd.n36 0.001
R906 pad.n138 pad.n131 4.52159
R907 pad.n486 pad.n485 4.52158
R908 pad.n484 pad.n458 4.5005
R909 pad.n477 pad.n476 4.5005
R910 pad.n469 pad.n29 4.5005
R911 pad.n498 pad.n497 4.5005
R912 pad.n28 pad.n24 4.5005
R913 pad.n450 pad.n21 4.5005
R914 pad.n449 pad.n18 4.5005
R915 pad.n448 pad.n15 4.5005
R916 pad.n37 pad.n12 4.5005
R917 pad.n440 pad.n9 4.5005
R918 pad.n439 pad.n6 4.5005
R919 pad.n438 pad.n3 4.5005
R920 pad.n421 pad.n43 4.5005
R921 pad.n430 pad.n429 4.5005
R922 pad.n312 pad.n49 4.5005
R923 pad.n300 pad.n80 4.5005
R924 pad.n377 pad.n376 4.5005
R925 pad.n79 pad.n75 4.5005
R926 pad.n367 pad.n72 4.5005
R927 pad.n366 pad.n68 4.5005
R928 pad.n365 pad.n65 4.5005
R929 pad.n348 pad.n88 4.5005
R930 pad.n357 pad.n356 4.5005
R931 pad.n98 pad.n94 4.5005
R932 pad.n212 pad.n211 4.5005
R933 pad.n195 pad.n103 4.5005
R934 pad.n203 pad.n202 4.5005
R935 pad.n113 pad.n109 4.5005
R936 pad.n175 pad.n174 4.5005
R937 pad.n158 pad.n118 4.5005
R938 pad.n166 pad.n165 4.5005
R939 pad.n128 pad.n124 4.5005
R940 pad.n137 pad.n136 4.5005
R941 pad.n132 pad.n131 4.5005
R942 pad.n136 pad.n135 4.5005
R943 pad.n124 pad.n123 4.5005
R944 pad.n167 pad.n166 4.5005
R945 pad.n119 pad.n118 4.5005
R946 pad.n174 pad.n173 4.5005
R947 pad.n109 pad.n108 4.5005
R948 pad.n204 pad.n203 4.5005
R949 pad.n104 pad.n103 4.5005
R950 pad.n211 pad.n210 4.5005
R951 pad.n94 pad.n93 4.5005
R952 pad.n358 pad.n357 4.5005
R953 pad.n89 pad.n88 4.5005
R954 pad.n365 pad.n364 4.5005
R955 pad.n366 pad.n87 4.5005
R956 pad.n368 pad.n367 4.5005
R957 pad.n81 pad.n79 4.5005
R958 pad.n376 pad.n375 4.5005
R959 pad.n82 pad.n80 4.5005
R960 pad.n49 pad.n48 4.5005
R961 pad.n431 pad.n430 4.5005
R962 pad.n44 pad.n43 4.5005
R963 pad.n438 pad.n437 4.5005
R964 pad.n439 pad.n42 4.5005
R965 pad.n441 pad.n440 4.5005
R966 pad.n38 pad.n37 4.5005
R967 pad.n448 pad.n447 4.5005
R968 pad.n449 pad.n36 4.5005
R969 pad.n451 pad.n450 4.5005
R970 pad.n30 pad.n28 4.5005
R971 pad.n497 pad.n496 4.5005
R972 pad.n31 pad.n29 4.5005
R973 pad.n476 pad.n456 4.5005
R974 pad.n458 pad.n457 4.5005
R975 pad.n487 pad.n486 4.5005
R976 pad.n248 pad.n53 4.47552
R977 pad.n319 pad.n290 4.47552
R978 pad.n324 pad.n323 4.47552
R979 pad.n275 pad.n274 4.47552
R980 pad.n332 pad.n329 4.47552
R981 pad.n282 pad.n62 4.47552
R982 pad.n337 pad.n227 4.47552
R983 pad.n264 pad.n262 4.47552
R984 pad.n253 pad.n252 3.07063
R985 pad.n233 pad.n227 3.07063
R986 pad.n337 pad.n336 3.07063
R987 pad.n338 pad.n56 3.07063
R988 pad.n277 pad.n276 3.0005
R989 pad.n268 pad.n239 3.0005
R990 pad.n288 pad.n287 3.0005
R991 pad.n250 pad.n249 3.0005
R992 pad.n279 pad.n230 3.0005
R993 pad.n329 pad.n328 3.0005
R994 pad.n275 pad.n232 3.0005
R995 pad.n325 pad.n324 3.0005
R996 pad.n290 pad.n289 3.0005
R997 pad.n248 pad.n247 3.0005
R998 pad.n282 pad.n281 3.0005
R999 pad.n284 pad.n283 3.0005
R1000 pad.n335 pad.n62 3.0005
R1001 pad.n333 pad.n332 3.0005
R1002 pad.n274 pad.n273 3.0005
R1003 pad.n323 pad.n322 3.0005
R1004 pad.n320 pad.n319 3.0005
R1005 pad.n258 pad.n53 3.0005
R1006 pad.n407 pad.n406 3.0005
R1007 pad.n331 pad.n61 3.0005
R1008 pad.n272 pad.n271 3.0005
R1009 pad.n241 pad.n240 3.0005
R1010 pad.n318 pad.n317 3.0005
R1011 pad.n411 pad.n410 3.0005
R1012 pad.n257 pad.n55 3.0005
R1013 pad.n262 pad.n261 3.0005
R1014 pad.n264 pad.n263 3.0005
R1015 pad.n266 pad.n265 3.0005
R1016 pad.n280 pad.t3 2.31826
R1017 pad.n229 pad.t0 2.31826
R1018 pad.n246 pad.t12 2.31826
R1019 pad.n244 pad.t10 2.31826
R1020 pad.n238 pad.t9 2.31826
R1021 pad.n269 pad.t7 2.31826
R1022 pad.n251 pad.t14 2.31791
R1023 pad.n256 pad.t4 2.31592
R1024 pad.n133 pad.n132 2.20699
R1025 pad.n489 pad.n487 2.2005
R1026 pad.n490 pad.n457 2.2005
R1027 pad.n491 pad.n456 2.2005
R1028 pad.n33 pad.n31 2.2005
R1029 pad.n496 pad.n495 2.2005
R1030 pad.n32 pad.n30 2.2005
R1031 pad.n452 pad.n451 2.2005
R1032 pad.n36 pad.n35 2.2005
R1033 pad.n447 pad.n446 2.2005
R1034 pad.n39 pad.n38 2.2005
R1035 pad.n442 pad.n441 2.2005
R1036 pad.n42 pad.n41 2.2005
R1037 pad.n437 pad.n436 2.2005
R1038 pad.n45 pad.n44 2.2005
R1039 pad.n432 pad.n431 2.2005
R1040 pad.n48 pad.n47 2.2005
R1041 pad.n84 pad.n82 2.2005
R1042 pad.n375 pad.n374 2.2005
R1043 pad.n83 pad.n81 2.2005
R1044 pad.n369 pad.n368 2.2005
R1045 pad.n87 pad.n86 2.2005
R1046 pad.n364 pad.n363 2.2005
R1047 pad.n90 pad.n89 2.2005
R1048 pad.n359 pad.n358 2.2005
R1049 pad.n93 pad.n92 2.2005
R1050 pad.n210 pad.n209 2.2005
R1051 pad.n105 pad.n104 2.2005
R1052 pad.n205 pad.n204 2.2005
R1053 pad.n108 pad.n107 2.2005
R1054 pad.n173 pad.n172 2.2005
R1055 pad.n120 pad.n119 2.2005
R1056 pad.n168 pad.n167 2.2005
R1057 pad.n123 pad.n122 2.2005
R1058 pad.n135 pad.n134 2.2005
R1059 pad.n412 pad.t19 1.78531
R1060 pad.n316 pad.t17 1.78531
R1061 pad.n295 pad.t22 1.78531
R1062 pad.n270 pad.t16 1.78531
R1063 pad.n330 pad.t18 1.78531
R1064 pad.n405 pad.t20 1.78531
R1065 pad.n0 pad.t21 1.78531
R1066 pad.n339 pad.t23 1.78502
R1067 pad.n483 pad.n459 1.5005
R1068 pad.n482 pad.n481 1.5005
R1069 pad.n480 pad.n460 1.5005
R1070 pad.n479 pad.n478 1.5005
R1071 pad.n475 pad.n461 1.5005
R1072 pad.n474 pad.n473 1.5005
R1073 pad.n472 pad.n462 1.5005
R1074 pad.n471 pad.n470 1.5005
R1075 pad.n468 pad.n463 1.5005
R1076 pad.n467 pad.n466 1.5005
R1077 pad.n465 pad.n464 1.5005
R1078 pad.n27 pad.n26 1.5005
R1079 pad.n500 pad.n499 1.5005
R1080 pad.n501 pad.n25 1.5005
R1081 pad.n503 pad.n502 1.5005
R1082 pad.n504 pad.n23 1.5005
R1083 pad.n506 pad.n505 1.5005
R1084 pad.n507 pad.n22 1.5005
R1085 pad.n509 pad.n508 1.5005
R1086 pad.n510 pad.n20 1.5005
R1087 pad.n512 pad.n511 1.5005
R1088 pad.n513 pad.n19 1.5005
R1089 pad.n515 pad.n514 1.5005
R1090 pad.n516 pad.n17 1.5005
R1091 pad.n518 pad.n517 1.5005
R1092 pad.n519 pad.n16 1.5005
R1093 pad.n521 pad.n520 1.5005
R1094 pad.n522 pad.n14 1.5005
R1095 pad.n524 pad.n523 1.5005
R1096 pad.n525 pad.n13 1.5005
R1097 pad.n527 pad.n526 1.5005
R1098 pad.n528 pad.n11 1.5005
R1099 pad.n530 pad.n529 1.5005
R1100 pad.n531 pad.n10 1.5005
R1101 pad.n533 pad.n532 1.5005
R1102 pad.n534 pad.n8 1.5005
R1103 pad.n536 pad.n535 1.5005
R1104 pad.n537 pad.n7 1.5005
R1105 pad.n539 pad.n538 1.5005
R1106 pad.n540 pad.n5 1.5005
R1107 pad.n542 pad.n541 1.5005
R1108 pad.n543 pad.n4 1.5005
R1109 pad.n545 pad.n544 1.5005
R1110 pad.n546 pad.n2 1.5005
R1111 pad.n548 pad.n547 1.5005
R1112 pad.n415 pad.n1 1.5005
R1113 pad.n417 pad.n416 1.5005
R1114 pad.n418 pad.n414 1.5005
R1115 pad.n420 pad.n419 1.5005
R1116 pad.n422 pad.n413 1.5005
R1117 pad.n424 pad.n423 1.5005
R1118 pad.n425 pad.n51 1.5005
R1119 pad.n428 pad.n427 1.5005
R1120 pad.n52 pad.n50 1.5005
R1121 pad.n308 pad.n307 1.5005
R1122 pad.n310 pad.n309 1.5005
R1123 pad.n311 pad.n292 1.5005
R1124 pad.n314 pad.n313 1.5005
R1125 pad.n306 pad.n291 1.5005
R1126 pad.n305 pad.n304 1.5005
R1127 pad.n303 pad.n293 1.5005
R1128 pad.n302 pad.n301 1.5005
R1129 pad.n299 pad.n294 1.5005
R1130 pad.n298 pad.n297 1.5005
R1131 pad.n78 pad.n77 1.5005
R1132 pad.n378 pad.n377 1.5005
R1133 pad.n379 pad.n76 1.5005
R1134 pad.n381 pad.n380 1.5005
R1135 pad.n382 pad.n74 1.5005
R1136 pad.n384 pad.n383 1.5005
R1137 pad.n386 pad.n73 1.5005
R1138 pad.n388 pad.n387 1.5005
R1139 pad.n389 pad.n71 1.5005
R1140 pad.n391 pad.n390 1.5005
R1141 pad.n392 pad.n69 1.5005
R1142 pad.n394 pad.n393 1.5005
R1143 pad.n395 pad.n67 1.5005
R1144 pad.n397 pad.n396 1.5005
R1145 pad.n398 pad.n66 1.5005
R1146 pad.n400 pad.n399 1.5005
R1147 pad.n401 pad.n64 1.5005
R1148 pad.n403 pad.n402 1.5005
R1149 pad.n342 pad.n63 1.5005
R1150 pad.n344 pad.n343 1.5005
R1151 pad.n345 pad.n341 1.5005
R1152 pad.n347 pad.n346 1.5005
R1153 pad.n349 pad.n340 1.5005
R1154 pad.n351 pad.n350 1.5005
R1155 pad.n352 pad.n96 1.5005
R1156 pad.n355 pad.n354 1.5005
R1157 pad.n226 pad.n95 1.5005
R1158 pad.n225 pad.n224 1.5005
R1159 pad.n223 pad.n97 1.5005
R1160 pad.n222 pad.n221 1.5005
R1161 pad.n220 pad.n219 1.5005
R1162 pad.n218 pad.n99 1.5005
R1163 pad.n217 pad.n216 1.5005
R1164 pad.n215 pad.n100 1.5005
R1165 pad.n214 pad.n213 1.5005
R1166 pad.n102 pad.n101 1.5005
R1167 pad.n192 pad.n191 1.5005
R1168 pad.n194 pad.n193 1.5005
R1169 pad.n196 pad.n190 1.5005
R1170 pad.n198 pad.n197 1.5005
R1171 pad.n199 pad.n111 1.5005
R1172 pad.n201 pad.n200 1.5005
R1173 pad.n189 pad.n110 1.5005
R1174 pad.n188 pad.n187 1.5005
R1175 pad.n186 pad.n112 1.5005
R1176 pad.n185 pad.n184 1.5005
R1177 pad.n183 pad.n182 1.5005
R1178 pad.n181 pad.n114 1.5005
R1179 pad.n180 pad.n179 1.5005
R1180 pad.n178 pad.n115 1.5005
R1181 pad.n177 pad.n176 1.5005
R1182 pad.n117 pad.n116 1.5005
R1183 pad.n154 pad.n153 1.5005
R1184 pad.n155 pad.n152 1.5005
R1185 pad.n157 pad.n156 1.5005
R1186 pad.n159 pad.n151 1.5005
R1187 pad.n161 pad.n160 1.5005
R1188 pad.n162 pad.n126 1.5005
R1189 pad.n164 pad.n163 1.5005
R1190 pad.n150 pad.n125 1.5005
R1191 pad.n149 pad.n148 1.5005
R1192 pad.n147 pad.n127 1.5005
R1193 pad.n146 pad.n145 1.5005
R1194 pad.n144 pad.n143 1.5005
R1195 pad.n142 pad.n129 1.5005
R1196 pad.n141 pad.n140 1.5005
R1197 pad.n139 pad.n130 1.5005
R1198 pad.n412 pad.n411 1.36955
R1199 pad.n318 pad.n316 1.36955
R1200 pad.n295 pad.n241 1.36955
R1201 pad.n272 pad.n270 1.36955
R1202 pad.n331 pad.n330 1.36955
R1203 pad.n406 pad.n405 1.36955
R1204 pad.n339 pad.n338 1.36955
R1205 pad.n257 pad.n0 1.36955
R1206 pad.n256 pad.t5 1.294
R1207 pad.n280 pad.t6 1.294
R1208 pad.n229 pad.t2 1.294
R1209 pad.n246 pad.t13 1.294
R1210 pad.n244 pad.t1 1.294
R1211 pad.n238 pad.t11 1.294
R1212 pad.n269 pad.t8 1.294
R1213 pad.n251 pad.t15 1.29365
R1214 pad.n122 pad.n121 1.1005
R1215 pad.n169 pad.n168 1.1005
R1216 pad.n170 pad.n120 1.1005
R1217 pad.n172 pad.n171 1.1005
R1218 pad.n107 pad.n106 1.1005
R1219 pad.n206 pad.n205 1.1005
R1220 pad.n207 pad.n105 1.1005
R1221 pad.n209 pad.n208 1.1005
R1222 pad.n92 pad.n91 1.1005
R1223 pad.n360 pad.n359 1.1005
R1224 pad.n361 pad.n90 1.1005
R1225 pad.n363 pad.n362 1.1005
R1226 pad.n86 pad.n85 1.1005
R1227 pad.n370 pad.n369 1.1005
R1228 pad.n371 pad.n83 1.1005
R1229 pad.n374 pad.n373 1.1005
R1230 pad.n372 pad.n84 1.1005
R1231 pad.n47 pad.n46 1.1005
R1232 pad.n433 pad.n432 1.1005
R1233 pad.n434 pad.n45 1.1005
R1234 pad.n436 pad.n435 1.1005
R1235 pad.n41 pad.n40 1.1005
R1236 pad.n443 pad.n442 1.1005
R1237 pad.n444 pad.n39 1.1005
R1238 pad.n446 pad.n445 1.1005
R1239 pad.n35 pad.n34 1.1005
R1240 pad.n453 pad.n452 1.1005
R1241 pad.n454 pad.n32 1.1005
R1242 pad.n495 pad.n494 1.1005
R1243 pad.n493 pad.n33 1.1005
R1244 pad.n492 pad.n491 1.1005
R1245 pad.n490 pad.n455 1.1005
R1246 pad.n489 pad.n488 1.1005
R1247 pad.n249 pad 1.09761
R1248 pad.n288 pad 1.09761
R1249 pad.n239 pad 1.09761
R1250 pad.n276 pad 1.09761
R1251 pad.n230 pad 1.09761
R1252 pad.n283 pad 1.09761
R1253 pad.n252 pad 1.09761
R1254 pad.n265 pad 1.09761
R1255 pad.n426 pad 0.83073
R1256 pad pad.n315 0.83073
R1257 pad.n296 pad 0.83073
R1258 pad.n385 pad 0.83073
R1259 pad pad.n70 0.83073
R1260 pad pad.n404 0.83073
R1261 pad.n353 pad 0.83073
R1262 pad pad.n549 0.83073
R1263 pad.n286 pad.t26 0.672378
R1264 pad.t25 pad.n237 0.672378
R1265 pad.n243 pad.t24 0.672378
R1266 pad.t27 pad.n54 0.672378
R1267 pad.n249 pad.n248 0.64968
R1268 pad.n411 pad.n53 0.64968
R1269 pad.n290 pad.n288 0.64968
R1270 pad.n319 pad.n318 0.64968
R1271 pad.n324 pad.n239 0.64968
R1272 pad.n323 pad.n241 0.64968
R1273 pad.n276 pad.n275 0.64968
R1274 pad.n274 pad.n272 0.64968
R1275 pad.n329 pad.n230 0.64968
R1276 pad.n332 pad.n331 0.64968
R1277 pad.n283 pad.n282 0.64968
R1278 pad.n406 pad.n62 0.64968
R1279 pad.n252 pad.n227 0.64968
R1280 pad.n338 pad.n337 0.64968
R1281 pad.n265 pad.n264 0.64968
R1282 pad.n262 pad.n257 0.64968
R1283 pad.t26 pad.n267 0.589365
R1284 pad.t26 pad.n245 0.589365
R1285 pad.t26 pad.n278 0.589365
R1286 pad.t26 pad.n254 0.589365
R1287 pad.t26 pad.n285 0.589365
R1288 pad.t25 pad.n236 0.589365
R1289 pad.t25 pad.n234 0.589365
R1290 pad.t25 pad.n326 0.589365
R1291 pad.n327 pad.t25 0.589365
R1292 pad.t25 pad.n231 0.589365
R1293 pad.n259 pad.t24 0.589365
R1294 pad.n321 pad.t24 0.589365
R1295 pad.n242 pad.t24 0.589365
R1296 pad.n228 pad.t24 0.589365
R1297 pad.n334 pad.t24 0.589365
R1298 pad.n409 pad.t27 0.589365
R1299 pad.t27 pad.n58 0.589365
R1300 pad.t27 pad.n60 0.589365
R1301 pad.t27 pad.n57 0.589365
R1302 pad.t27 pad.n408 0.589365
R1303 pad.n133 pad.n121 0.557177
R1304 pad pad.n246 0.435451
R1305 pad pad.n244 0.435451
R1306 pad pad.n238 0.435451
R1307 pad pad.n269 0.435451
R1308 pad pad.n229 0.435451
R1309 pad pad.n280 0.435451
R1310 pad pad.n251 0.435451
R1311 pad pad.n256 0.435451
R1312 pad.t26 pad.n255 0.419935
R1313 pad.t25 pad.n235 0.419935
R1314 pad.n260 pad.t24 0.419935
R1315 pad.t27 pad.n59 0.419935
R1316 pad.t26 pad.n253 0.32731
R1317 pad.t25 pad.n233 0.32731
R1318 pad.n336 pad.t24 0.32731
R1319 pad.t27 pad.n56 0.32731
R1320 pad pad.n412 0.317156
R1321 pad.n316 pad 0.317156
R1322 pad pad.n295 0.317156
R1323 pad.n270 pad 0.317156
R1324 pad.n330 pad 0.317156
R1325 pad.n405 pad 0.317156
R1326 pad pad.n339 0.317156
R1327 pad pad.n0 0.317156
R1328 pad.n139 pad.n138 0.278474
R1329 pad.n485 pad.n459 0.278376
R1330 pad.n255 pad 0.188225
R1331 pad.n235 pad 0.188225
R1332 pad.n260 pad 0.188225
R1333 pad.n59 pad 0.188225
R1334 pad.n284 pad.n253 0.183954
R1335 pad.n281 pad.n233 0.183954
R1336 pad.n336 pad.n335 0.183954
R1337 pad.n407 pad.n56 0.183954
R1338 pad.n266 pad.n255 0.160165
R1339 pad.n263 pad.n235 0.160165
R1340 pad.n261 pad.n260 0.160165
R1341 pad.n59 pad.n55 0.160165
R1342 pad.n267 pad.n266 0.146012
R1343 pad.n263 pad.n236 0.146012
R1344 pad.n261 pad.n259 0.146012
R1345 pad.n409 pad.n55 0.146012
R1346 pad.n268 pad.n245 0.140121
R1347 pad.n325 pad.n234 0.140121
R1348 pad.n322 pad.n321 0.140121
R1349 pad.n240 pad.n58 0.140121
R1350 pad.n278 pad.n277 0.136629
R1351 pad.n326 pad.n232 0.136629
R1352 pad.n273 pad.n242 0.136629
R1353 pad.n271 pad.n60 0.136629
R1354 pad.n286 pad.n250 0.135252
R1355 pad.n247 pad.n237 0.135252
R1356 pad.n258 pad.n243 0.135252
R1357 pad.n410 pad.n54 0.135252
R1358 pad.n285 pad.n279 0.13379
R1359 pad.n328 pad.n231 0.13379
R1360 pad.n334 pad.n333 0.13379
R1361 pad.n408 pad.n61 0.13379
R1362 pad.n279 pad.n254 0.133137
R1363 pad.n328 pad.n327 0.133137
R1364 pad.n333 pad.n228 0.133137
R1365 pad.n61 pad.n57 0.133137
R1366 pad.n277 pad.n254 0.130298
R1367 pad.n327 pad.n232 0.130298
R1368 pad.n273 pad.n228 0.130298
R1369 pad.n271 pad.n57 0.130298
R1370 pad.n287 pad.n286 0.129894
R1371 pad.n289 pad.n237 0.129894
R1372 pad.n320 pad.n243 0.129894
R1373 pad.n317 pad.n54 0.129894
R1374 pad.n285 pad.n284 0.129645
R1375 pad.n281 pad.n231 0.129645
R1376 pad.n335 pad.n334 0.129645
R1377 pad.n408 pad.n407 0.129645
R1378 pad.n278 pad.n268 0.126806
R1379 pad.n326 pad.n325 0.126806
R1380 pad.n322 pad.n242 0.126806
R1381 pad.n240 pad.n60 0.126806
R1382 pad.n287 pad.n245 0.123314
R1383 pad.n289 pad.n234 0.123314
R1384 pad.n321 pad.n320 0.123314
R1385 pad.n317 pad.n58 0.123314
R1386 pad.n267 pad.n250 0.117423
R1387 pad.n247 pad.n236 0.117423
R1388 pad.n259 pad.n258 0.117423
R1389 pad.n410 pad.n409 0.117423
R1390 pad.n136 pad.n131 0.0591667
R1391 pad.n136 pad.n124 0.0591667
R1392 pad.n166 pad.n124 0.0591667
R1393 pad.n166 pad.n118 0.0591667
R1394 pad.n174 pad.n118 0.0591667
R1395 pad.n174 pad.n109 0.0591667
R1396 pad.n203 pad.n109 0.0591667
R1397 pad.n203 pad.n103 0.0591667
R1398 pad.n211 pad.n103 0.0591667
R1399 pad.n211 pad.n94 0.0591667
R1400 pad.n357 pad.n94 0.0591667
R1401 pad.n357 pad.n88 0.0591667
R1402 pad.n365 pad.n88 0.0591667
R1403 pad.n366 pad.n365 0.0591667
R1404 pad.n367 pad.n366 0.0591667
R1405 pad.n367 pad.n79 0.0591667
R1406 pad.n376 pad.n79 0.0591667
R1407 pad.n376 pad.n80 0.0591667
R1408 pad.n80 pad.n49 0.0591667
R1409 pad.n430 pad.n49 0.0591667
R1410 pad.n430 pad.n43 0.0591667
R1411 pad.n438 pad.n43 0.0591667
R1412 pad.n439 pad.n438 0.0591667
R1413 pad.n440 pad.n439 0.0591667
R1414 pad.n440 pad.n37 0.0591667
R1415 pad.n448 pad.n37 0.0591667
R1416 pad.n449 pad.n448 0.0591667
R1417 pad.n450 pad.n449 0.0591667
R1418 pad.n450 pad.n28 0.0591667
R1419 pad.n497 pad.n28 0.0591667
R1420 pad.n497 pad.n29 0.0591667
R1421 pad.n476 pad.n29 0.0591667
R1422 pad.n476 pad.n458 0.0591667
R1423 pad.n486 pad.n458 0.0591667
R1424 pad.n135 pad.n132 0.0591667
R1425 pad.n135 pad.n123 0.0591667
R1426 pad.n167 pad.n123 0.0591667
R1427 pad.n167 pad.n119 0.0591667
R1428 pad.n173 pad.n119 0.0591667
R1429 pad.n173 pad.n108 0.0591667
R1430 pad.n204 pad.n108 0.0591667
R1431 pad.n204 pad.n104 0.0591667
R1432 pad.n210 pad.n104 0.0591667
R1433 pad.n210 pad.n93 0.0591667
R1434 pad.n358 pad.n93 0.0591667
R1435 pad.n358 pad.n89 0.0591667
R1436 pad.n364 pad.n89 0.0591667
R1437 pad.n364 pad.n87 0.0591667
R1438 pad.n368 pad.n87 0.0591667
R1439 pad.n368 pad.n81 0.0591667
R1440 pad.n375 pad.n81 0.0591667
R1441 pad.n375 pad.n82 0.0591667
R1442 pad.n82 pad.n48 0.0591667
R1443 pad.n431 pad.n48 0.0591667
R1444 pad.n431 pad.n44 0.0591667
R1445 pad.n437 pad.n44 0.0591667
R1446 pad.n437 pad.n42 0.0591667
R1447 pad.n441 pad.n42 0.0591667
R1448 pad.n441 pad.n38 0.0591667
R1449 pad.n447 pad.n38 0.0591667
R1450 pad.n447 pad.n36 0.0591667
R1451 pad.n451 pad.n36 0.0591667
R1452 pad.n451 pad.n30 0.0591667
R1453 pad.n496 pad.n30 0.0591667
R1454 pad.n496 pad.n31 0.0591667
R1455 pad.n456 pad.n31 0.0591667
R1456 pad.n457 pad.n456 0.0591667
R1457 pad.n487 pad.n457 0.0591667
R1458 pad.n485 pad.n484 0.0407494
R1459 pad.n138 pad.n137 0.0407425
R1460 pad.n140 pad.n139 0.0148733
R1461 pad.n140 pad.n129 0.0148733
R1462 pad.n144 pad.n129 0.0148733
R1463 pad.n145 pad.n144 0.0148733
R1464 pad.n145 pad.n127 0.0148733
R1465 pad.n149 pad.n127 0.0148733
R1466 pad.n150 pad.n149 0.0148733
R1467 pad.n163 pad.n150 0.0148733
R1468 pad.n163 pad.n162 0.0148733
R1469 pad.n162 pad.n161 0.0148733
R1470 pad.n161 pad.n151 0.0148733
R1471 pad.n156 pad.n151 0.0148733
R1472 pad.n156 pad.n155 0.0148733
R1473 pad.n155 pad.n154 0.0148733
R1474 pad.n154 pad.n116 0.0148733
R1475 pad.n177 pad.n116 0.0148733
R1476 pad.n178 pad.n177 0.0148733
R1477 pad.n179 pad.n178 0.0148733
R1478 pad.n179 pad.n114 0.0148733
R1479 pad.n183 pad.n114 0.0148733
R1480 pad.n184 pad.n183 0.0148733
R1481 pad.n184 pad.n112 0.0148733
R1482 pad.n188 pad.n112 0.0148733
R1483 pad.n189 pad.n188 0.0148733
R1484 pad.n200 pad.n189 0.0148733
R1485 pad.n200 pad.n199 0.0148733
R1486 pad.n199 pad.n198 0.0148733
R1487 pad.n198 pad.n190 0.0148733
R1488 pad.n193 pad.n190 0.0148733
R1489 pad.n193 pad.n192 0.0148733
R1490 pad.n192 pad.n101 0.0148733
R1491 pad.n214 pad.n101 0.0148733
R1492 pad.n215 pad.n214 0.0148733
R1493 pad.n216 pad.n215 0.0148733
R1494 pad.n216 pad.n99 0.0148733
R1495 pad.n220 pad.n99 0.0148733
R1496 pad.n221 pad.n220 0.0148733
R1497 pad.n221 pad.n97 0.0148733
R1498 pad.n225 pad.n97 0.0148733
R1499 pad.n226 pad.n225 0.0148733
R1500 pad.n354 pad.n226 0.0148733
R1501 pad.n352 pad.n351 0.0148733
R1502 pad.n351 pad.n340 0.0148733
R1503 pad.n346 pad.n340 0.0148733
R1504 pad.n346 pad.n345 0.0148733
R1505 pad.n345 pad.n344 0.0148733
R1506 pad.n344 pad.n63 0.0148733
R1507 pad.n403 pad.n64 0.0148733
R1508 pad.n399 pad.n64 0.0148733
R1509 pad.n399 pad.n398 0.0148733
R1510 pad.n398 pad.n397 0.0148733
R1511 pad.n397 pad.n67 0.0148733
R1512 pad.n393 pad.n392 0.0148733
R1513 pad.n392 pad.n391 0.0148733
R1514 pad.n391 pad.n71 0.0148733
R1515 pad.n387 pad.n71 0.0148733
R1516 pad.n387 pad.n386 0.0148733
R1517 pad.n384 pad.n74 0.0148733
R1518 pad.n380 pad.n74 0.0148733
R1519 pad.n380 pad.n379 0.0148733
R1520 pad.n379 pad.n378 0.0148733
R1521 pad.n378 pad.n77 0.0148733
R1522 pad.n297 pad.n294 0.0148733
R1523 pad.n302 pad.n294 0.0148733
R1524 pad.n303 pad.n302 0.0148733
R1525 pad.n304 pad.n303 0.0148733
R1526 pad.n304 pad.n291 0.0148733
R1527 pad.n314 pad.n292 0.0148733
R1528 pad.n309 pad.n292 0.0148733
R1529 pad.n309 pad.n308 0.0148733
R1530 pad.n308 pad.n52 0.0148733
R1531 pad.n427 pad.n52 0.0148733
R1532 pad.n425 pad.n424 0.0148733
R1533 pad.n424 pad.n413 0.0148733
R1534 pad.n419 pad.n413 0.0148733
R1535 pad.n419 pad.n418 0.0148733
R1536 pad.n418 pad.n417 0.0148733
R1537 pad.n417 pad.n1 0.0148733
R1538 pad.n548 pad.n2 0.0148733
R1539 pad.n544 pad.n2 0.0148733
R1540 pad.n544 pad.n543 0.0148733
R1541 pad.n543 pad.n542 0.0148733
R1542 pad.n542 pad.n5 0.0148733
R1543 pad.n538 pad.n5 0.0148733
R1544 pad.n538 pad.n537 0.0148733
R1545 pad.n537 pad.n536 0.0148733
R1546 pad.n536 pad.n8 0.0148733
R1547 pad.n532 pad.n8 0.0148733
R1548 pad.n532 pad.n531 0.0148733
R1549 pad.n531 pad.n530 0.0148733
R1550 pad.n530 pad.n11 0.0148733
R1551 pad.n526 pad.n11 0.0148733
R1552 pad.n526 pad.n525 0.0148733
R1553 pad.n525 pad.n524 0.0148733
R1554 pad.n524 pad.n14 0.0148733
R1555 pad.n520 pad.n14 0.0148733
R1556 pad.n520 pad.n519 0.0148733
R1557 pad.n519 pad.n518 0.0148733
R1558 pad.n518 pad.n17 0.0148733
R1559 pad.n514 pad.n17 0.0148733
R1560 pad.n514 pad.n513 0.0148733
R1561 pad.n513 pad.n512 0.0148733
R1562 pad.n512 pad.n20 0.0148733
R1563 pad.n508 pad.n20 0.0148733
R1564 pad.n508 pad.n507 0.0148733
R1565 pad.n507 pad.n506 0.0148733
R1566 pad.n506 pad.n23 0.0148733
R1567 pad.n502 pad.n23 0.0148733
R1568 pad.n502 pad.n501 0.0148733
R1569 pad.n501 pad.n500 0.0148733
R1570 pad.n500 pad.n26 0.0148733
R1571 pad.n465 pad.n26 0.0148733
R1572 pad.n466 pad.n465 0.0148733
R1573 pad.n466 pad.n463 0.0148733
R1574 pad.n471 pad.n463 0.0148733
R1575 pad.n472 pad.n471 0.0148733
R1576 pad.n473 pad.n472 0.0148733
R1577 pad.n473 pad.n461 0.0148733
R1578 pad.n479 pad.n461 0.0148733
R1579 pad.n480 pad.n479 0.0148733
R1580 pad.n481 pad.n480 0.0148733
R1581 pad.n481 pad.n459 0.0148733
R1582 pad.n141 pad.n130 0.0148733
R1583 pad.n142 pad.n141 0.0148733
R1584 pad.n143 pad.n142 0.0148733
R1585 pad.n147 pad.n146 0.0148733
R1586 pad.n148 pad.n147 0.0148733
R1587 pad.n148 pad.n125 0.0148733
R1588 pad.n164 pad.n126 0.0148733
R1589 pad.n160 pad.n126 0.0148733
R1590 pad.n160 pad.n159 0.0148733
R1591 pad.n157 pad.n152 0.0148733
R1592 pad.n153 pad.n152 0.0148733
R1593 pad.n153 pad.n117 0.0148733
R1594 pad.n176 pad.n117 0.0148733
R1595 pad.n180 pad.n115 0.0148733
R1596 pad.n181 pad.n180 0.0148733
R1597 pad.n182 pad.n181 0.0148733
R1598 pad.n186 pad.n185 0.0148733
R1599 pad.n187 pad.n186 0.0148733
R1600 pad.n187 pad.n110 0.0148733
R1601 pad.n201 pad.n111 0.0148733
R1602 pad.n197 pad.n111 0.0148733
R1603 pad.n197 pad.n196 0.0148733
R1604 pad.n194 pad.n191 0.0148733
R1605 pad.n191 pad.n102 0.0148733
R1606 pad.n213 pad.n102 0.0148733
R1607 pad.n217 pad.n100 0.0148733
R1608 pad.n218 pad.n217 0.0148733
R1609 pad.n219 pad.n218 0.0148733
R1610 pad.n223 pad.n222 0.0148733
R1611 pad.n224 pad.n223 0.0148733
R1612 pad.n224 pad.n95 0.0148733
R1613 pad.n355 pad.n96 0.0148733
R1614 pad.n350 pad.n96 0.0148733
R1615 pad.n350 pad.n349 0.0148733
R1616 pad.n347 pad.n341 0.0148733
R1617 pad.n343 pad.n341 0.0148733
R1618 pad.n343 pad.n342 0.0148733
R1619 pad.n402 pad.n401 0.0148733
R1620 pad.n401 pad.n400 0.0148733
R1621 pad.n400 pad.n66 0.0148733
R1622 pad.n396 pad.n395 0.0148733
R1623 pad.n395 pad.n394 0.0148733
R1624 pad.n394 pad.n69 0.0148733
R1625 pad.n390 pad.n389 0.0148733
R1626 pad.n389 pad.n388 0.0148733
R1627 pad.n388 pad.n73 0.0148733
R1628 pad.n383 pad.n382 0.0148733
R1629 pad.n382 pad.n381 0.0148733
R1630 pad.n381 pad.n76 0.0148733
R1631 pad.n377 pad.n76 0.0148733
R1632 pad.n377 pad.n78 0.0148733
R1633 pad.n298 pad.n78 0.0148733
R1634 pad.n299 pad.n298 0.0148733
R1635 pad.n301 pad.n299 0.0148733
R1636 pad.n305 pad.n293 0.0148733
R1637 pad.n306 pad.n305 0.0148733
R1638 pad.n313 pad.n306 0.0148733
R1639 pad.n311 pad.n310 0.0148733
R1640 pad.n310 pad.n307 0.0148733
R1641 pad.n307 pad.n50 0.0148733
R1642 pad.n428 pad.n51 0.0148733
R1643 pad.n423 pad.n51 0.0148733
R1644 pad.n423 pad.n422 0.0148733
R1645 pad.n420 pad.n414 0.0148733
R1646 pad.n416 pad.n414 0.0148733
R1647 pad.n416 pad.n415 0.0148733
R1648 pad.n547 pad.n546 0.0148733
R1649 pad.n546 pad.n545 0.0148733
R1650 pad.n545 pad.n4 0.0148733
R1651 pad.n541 pad.n540 0.0148733
R1652 pad.n540 pad.n539 0.0148733
R1653 pad.n539 pad.n7 0.0148733
R1654 pad.n535 pad.n534 0.0148733
R1655 pad.n534 pad.n533 0.0148733
R1656 pad.n533 pad.n10 0.0148733
R1657 pad.n529 pad.n528 0.0148733
R1658 pad.n528 pad.n527 0.0148733
R1659 pad.n527 pad.n13 0.0148733
R1660 pad.n523 pad.n522 0.0148733
R1661 pad.n522 pad.n521 0.0148733
R1662 pad.n521 pad.n16 0.0148733
R1663 pad.n517 pad.n516 0.0148733
R1664 pad.n516 pad.n515 0.0148733
R1665 pad.n515 pad.n19 0.0148733
R1666 pad.n511 pad.n510 0.0148733
R1667 pad.n510 pad.n509 0.0148733
R1668 pad.n509 pad.n22 0.0148733
R1669 pad.n505 pad.n504 0.0148733
R1670 pad.n504 pad.n503 0.0148733
R1671 pad.n503 pad.n25 0.0148733
R1672 pad.n499 pad.n25 0.0148733
R1673 pad.n464 pad.n27 0.0148733
R1674 pad.n467 pad.n464 0.0148733
R1675 pad.n468 pad.n467 0.0148733
R1676 pad.n470 pad.n462 0.0148733
R1677 pad.n474 pad.n462 0.0148733
R1678 pad.n475 pad.n474 0.0148733
R1679 pad.n478 pad.n460 0.0148733
R1680 pad.n482 pad.n460 0.0148733
R1681 pad.n483 pad.n482 0.0148733
R1682 pad.n175 pad.n115 0.01458
R1683 pad.n24 pad.n22 0.01458
R1684 pad.n549 pad.n548 0.0144333
R1685 pad.n404 pad.n403 0.01414
R1686 pad.n159 pad.n158 0.0139933
R1687 pad.n498 pad.n27 0.0139933
R1688 pad.n75 pad.n73 0.0137
R1689 pad.n300 pad.n293 0.0137
R1690 pad.n185 pad.n113 0.0134067
R1691 pad.n21 pad.n19 0.0134067
R1692 pad.n354 pad.n353 0.01326
R1693 pad.n427 pad.n426 0.0129667
R1694 pad.n165 pad.n125 0.01282
R1695 pad.n470 pad.n469 0.01282
R1696 pad.n72 pad.n69 0.0125267
R1697 pad.n312 pad.n311 0.0125267
R1698 pad.n134 pad.n122 0.0125
R1699 pad.n168 pad.n122 0.0125
R1700 pad.n168 pad.n120 0.0125
R1701 pad.n172 pad.n120 0.0125
R1702 pad.n172 pad.n107 0.0125
R1703 pad.n205 pad.n107 0.0125
R1704 pad.n205 pad.n105 0.0125
R1705 pad.n209 pad.n105 0.0125
R1706 pad.n209 pad.n92 0.0125
R1707 pad.n359 pad.n92 0.0125
R1708 pad.n359 pad.n90 0.0125
R1709 pad.n363 pad.n90 0.0125
R1710 pad.n363 pad.n86 0.0125
R1711 pad.n369 pad.n86 0.0125
R1712 pad.n369 pad.n83 0.0125
R1713 pad.n374 pad.n83 0.0125
R1714 pad.n374 pad.n84 0.0125
R1715 pad.n84 pad.n47 0.0125
R1716 pad.n432 pad.n47 0.0125
R1717 pad.n432 pad.n45 0.0125
R1718 pad.n436 pad.n45 0.0125
R1719 pad.n436 pad.n41 0.0125
R1720 pad.n442 pad.n41 0.0125
R1721 pad.n442 pad.n39 0.0125
R1722 pad.n446 pad.n39 0.0125
R1723 pad.n446 pad.n35 0.0125
R1724 pad.n452 pad.n35 0.0125
R1725 pad.n452 pad.n32 0.0125
R1726 pad.n495 pad.n32 0.0125
R1727 pad.n495 pad.n33 0.0125
R1728 pad.n491 pad.n33 0.0125
R1729 pad.n491 pad.n490 0.0125
R1730 pad.n490 pad.n489 0.0125
R1731 pad.n202 pad.n201 0.0122333
R1732 pad.n18 pad.n16 0.0122333
R1733 pad.n393 pad.n70 0.0117933
R1734 pad.n143 pad.n128 0.0116467
R1735 pad.n478 pad.n477 0.0116467
R1736 pad.n68 pad.n66 0.0113533
R1737 pad.n429 pad.n428 0.0113533
R1738 pad.n195 pad.n194 0.01106
R1739 pad.n15 pad.n13 0.01106
R1740 pad.n315 pad.n291 0.01062
R1741 pad.n342 pad.n65 0.01018
R1742 pad.n421 pad.n420 0.01018
R1743 pad.n212 pad.n100 0.00988667
R1744 pad.n12 pad.n10 0.00988667
R1745 pad.n385 pad.n384 0.00944667
R1746 pad.n349 pad.n348 0.00900667
R1747 pad.n547 pad.n3 0.00900667
R1748 pad.n222 pad.n98 0.00871333
R1749 pad.n9 pad.n7 0.00871333
R1750 pad.n296 pad.n77 0.00827333
R1751 pad.n356 pad.n95 0.00783333
R1752 pad.n541 pad.n6 0.00783333
R1753 pad.n169 pad.n121 0.00783333
R1754 pad.n170 pad.n169 0.00783333
R1755 pad.n171 pad.n170 0.00783333
R1756 pad.n171 pad.n106 0.00783333
R1757 pad.n206 pad.n106 0.00783333
R1758 pad.n207 pad.n206 0.00783333
R1759 pad.n208 pad.n207 0.00783333
R1760 pad.n208 pad.n91 0.00783333
R1761 pad.n360 pad.n91 0.00783333
R1762 pad.n361 pad.n360 0.00783333
R1763 pad.n362 pad.n361 0.00783333
R1764 pad.n362 pad.n85 0.00783333
R1765 pad.n370 pad.n85 0.00783333
R1766 pad.n371 pad.n370 0.00783333
R1767 pad.n373 pad.n371 0.00783333
R1768 pad.n373 pad.n372 0.00783333
R1769 pad.n372 pad.n46 0.00783333
R1770 pad.n433 pad.n46 0.00783333
R1771 pad.n434 pad.n433 0.00783333
R1772 pad.n435 pad.n434 0.00783333
R1773 pad.n435 pad.n40 0.00783333
R1774 pad.n443 pad.n40 0.00783333
R1775 pad.n444 pad.n443 0.00783333
R1776 pad.n445 pad.n444 0.00783333
R1777 pad.n445 pad.n34 0.00783333
R1778 pad.n453 pad.n34 0.00783333
R1779 pad.n454 pad.n453 0.00783333
R1780 pad.n494 pad.n454 0.00783333
R1781 pad.n494 pad.n493 0.00783333
R1782 pad.n493 pad.n492 0.00783333
R1783 pad.n492 pad.n455 0.00783333
R1784 pad.n488 pad.n455 0.00783333
R1785 pad.n356 pad.n355 0.00754
R1786 pad.n6 pad.n4 0.00754
R1787 pad.n297 pad.n296 0.0071
R1788 pad.n134 pad.n133 0.00694773
R1789 pad.n219 pad.n98 0.00666
R1790 pad.n535 pad.n9 0.00666
R1791 pad.n348 pad.n347 0.00636667
R1792 pad.n415 pad.n3 0.00636667
R1793 pad.n386 pad.n385 0.00592667
R1794 pad.n213 pad.n212 0.00548667
R1795 pad.n529 pad.n12 0.00548667
R1796 pad.n402 pad.n65 0.00519333
R1797 pad.n422 pad.n421 0.00519333
R1798 pad.n137 pad.n130 0.0049
R1799 pad.n484 pad.n483 0.0049
R1800 pad.n315 pad.n314 0.00475333
R1801 pad.n196 pad.n195 0.00431333
R1802 pad.n523 pad.n15 0.00431333
R1803 pad.n488 pad 0.00416667
R1804 pad.n396 pad.n68 0.00402
R1805 pad.n429 pad.n50 0.00402
R1806 pad.n146 pad.n128 0.00372667
R1807 pad.n477 pad.n475 0.00372667
R1808 pad.n70 pad.n67 0.00358
R1809 pad.n202 pad.n110 0.00314
R1810 pad.n517 pad.n18 0.00314
R1811 pad.n390 pad.n72 0.00284667
R1812 pad.n313 pad.n312 0.00284667
R1813 pad.n165 pad.n164 0.00255333
R1814 pad.n469 pad.n468 0.00255333
R1815 pad.n426 pad.n425 0.00240667
R1816 pad.n353 pad.n352 0.00211333
R1817 pad.n182 pad.n113 0.00196667
R1818 pad.n511 pad.n21 0.00196667
R1819 pad.n383 pad.n75 0.00167333
R1820 pad.n301 pad.n300 0.00167333
R1821 pad.n158 pad.n157 0.00138
R1822 pad.n499 pad.n498 0.00138
R1823 pad.n404 pad.n63 0.00123333
R1824 pad.n549 pad.n1 0.00094
R1825 pad.n176 pad.n175 0.000793333
R1826 pad.n505 pad.n24 0.000793333
R1827 sg13g2_GateDecode_0.sg13g2_LevelUp_0.o sg13g2_Clamp_N15N15D_0.gate 66.1076
R1828 sg13g2_GateDecode_0.ngate.t0 sg13g2_GateDecode_0.ngate.n0 17.0005
R1829 sg13g2_GateDecode_0.ngate.n16 sg13g2_GateDecode_0.ngate.n15 9.75711
R1830 sg13g2_GateDecode_0.ngate.n2 sg13g2_GateDecode_0.ngate.t3 9.10182
R1831 sg13g2_GateDecode_0.ngate.n14 sg13g2_GateDecode_0.ngate.t2 8.24932
R1832 sg13g2_GateDecode_0.ngate.n13 sg13g2_GateDecode_0.ngate.t7 8.24932
R1833 sg13g2_GateDecode_0.ngate.n12 sg13g2_GateDecode_0.ngate.t13 8.24932
R1834 sg13g2_GateDecode_0.ngate.n11 sg13g2_GateDecode_0.ngate.t4 8.24932
R1835 sg13g2_GateDecode_0.ngate.n10 sg13g2_GateDecode_0.ngate.t14 8.24932
R1836 sg13g2_GateDecode_0.ngate.n9 sg13g2_GateDecode_0.ngate.t17 8.24932
R1837 sg13g2_GateDecode_0.ngate.n8 sg13g2_GateDecode_0.ngate.t6 8.24932
R1838 sg13g2_GateDecode_0.ngate.n7 sg13g2_GateDecode_0.ngate.t16 8.24932
R1839 sg13g2_GateDecode_0.ngate.n6 sg13g2_GateDecode_0.ngate.t8 8.24932
R1840 sg13g2_GateDecode_0.ngate.n5 sg13g2_GateDecode_0.ngate.t9 8.24932
R1841 sg13g2_GateDecode_0.ngate.n4 sg13g2_GateDecode_0.ngate.t5 8.24932
R1842 sg13g2_GateDecode_0.ngate.n3 sg13g2_GateDecode_0.ngate.t11 8.24932
R1843 sg13g2_GateDecode_0.ngate.n2 sg13g2_GateDecode_0.ngate.t15 8.24932
R1844 sg13g2_GateDecode_0.ngate.n15 sg13g2_GateDecode_0.ngate.t10 8.24932
R1845 sg13g2_GateDecode_0.ngate.n0 sg13g2_GateDecode_0.ngate.t1 4.53355
R1846 sg13g2_GateDecode_0.ngate.n17 sg13g2_GateDecode_0.ngate.n16 4.5005
R1847 sg13g2_GateDecode_0.ngate.n16 sg13g2_GateDecode_0.ngate.t12 4.31293
R1848 sg13g2_GateDecode_0.ngate.n1 sg13g2_GateDecode_0.ngate.t0 2.28308
R1849 sg13g2_GateDecode_0.sg13g2_LevelUp_0.o sg13g2_GateDecode_0.ngate.n1 1.9798
R1850 sg13g2_GateDecode_0.ngate.n3 sg13g2_GateDecode_0.ngate.n2 1.22425
R1851 sg13g2_GateDecode_0.ngate.n5 sg13g2_GateDecode_0.ngate.n4 1.22425
R1852 sg13g2_GateDecode_0.ngate.n7 sg13g2_GateDecode_0.ngate.n6 1.22425
R1853 sg13g2_GateDecode_0.ngate.n9 sg13g2_GateDecode_0.ngate.n8 1.22425
R1854 sg13g2_GateDecode_0.ngate.n11 sg13g2_GateDecode_0.ngate.n10 1.22425
R1855 sg13g2_GateDecode_0.ngate.n13 sg13g2_GateDecode_0.ngate.n12 1.22425
R1856 sg13g2_GateDecode_0.ngate.n15 sg13g2_GateDecode_0.ngate.n14 1.22425
R1857 sg13g2_Clamp_N15N15D_0.gate sg13g2_GateDecode_0.ngate.n17 1.17264
R1858 sg13g2_GateDecode_0.ngate.n4 sg13g2_GateDecode_0.ngate.n3 0.853
R1859 sg13g2_GateDecode_0.ngate.n6 sg13g2_GateDecode_0.ngate.n5 0.853
R1860 sg13g2_GateDecode_0.ngate.n8 sg13g2_GateDecode_0.ngate.n7 0.853
R1861 sg13g2_GateDecode_0.ngate.n10 sg13g2_GateDecode_0.ngate.n9 0.853
R1862 sg13g2_GateDecode_0.ngate.n12 sg13g2_GateDecode_0.ngate.n11 0.853
R1863 sg13g2_GateDecode_0.ngate.n14 sg13g2_GateDecode_0.ngate.n13 0.853
R1864 sg13g2_GateDecode_0.ngate.n17 sg13g2_Clamp_N15N15D_0.gate 0.1545
R1865 sg13g2_GateDecode_0.ngate.n1 sg13g2_GateDecode_0.ngate.n0 0.0738333
R1866 iovss.n220 iovss.n219 0.826084
R1867 iovss.n84 iovss.n80 0.826084
R1868 iovss.n218 iovss.n217 0.818682
R1869 iovss.n5 iovss.n4 0.818682
R1870 iovss.n206 iovss.n205 0.818682
R1871 iovss.n204 iovss.n12 0.818682
R1872 iovss.n203 iovss.n202 0.818682
R1873 iovss.n14 iovss.n13 0.818682
R1874 iovss.n191 iovss.n190 0.818682
R1875 iovss.n189 iovss.n21 0.818682
R1876 iovss.n188 iovss.n187 0.818682
R1877 iovss.n23 iovss.n22 0.818682
R1878 iovss.n176 iovss.n175 0.818682
R1879 iovss.n174 iovss.n30 0.818682
R1880 iovss.n173 iovss.n172 0.818682
R1881 iovss.n32 iovss.n31 0.818682
R1882 iovss.n161 iovss.n160 0.818682
R1883 iovss.n159 iovss.n39 0.818682
R1884 iovss.n158 iovss.n157 0.818682
R1885 iovss.n41 iovss.n40 0.818682
R1886 iovss.n146 iovss.n145 0.818682
R1887 iovss.n144 iovss.n48 0.818682
R1888 iovss.n143 iovss.n142 0.818682
R1889 iovss.n50 iovss.n49 0.818682
R1890 iovss.n131 iovss.n130 0.818682
R1891 iovss.n129 iovss.n57 0.818682
R1892 iovss.n128 iovss.n127 0.818682
R1893 iovss.n59 iovss.n58 0.818682
R1894 iovss.n116 iovss.n115 0.818682
R1895 iovss.n114 iovss.n66 0.818682
R1896 iovss.n113 iovss.n112 0.818682
R1897 iovss.n68 iovss.n67 0.818682
R1898 iovss.n101 iovss.n100 0.818682
R1899 iovss.n99 iovss.n75 0.818682
R1900 iovss.n98 iovss.n97 0.818682
R1901 iovss.n77 iovss.n76 0.818682
R1902 iovss.n86 iovss.n85 0.818682
R1903 iovss.n83 iovss.n81 0.818682
R1904 iovss.n87 iovss.n86 0.818682
R1905 iovss.n78 iovss.n77 0.818682
R1906 iovss.n97 iovss.n96 0.818682
R1907 iovss.n75 iovss.n73 0.818682
R1908 iovss.n102 iovss.n101 0.818682
R1909 iovss.n69 iovss.n68 0.818682
R1910 iovss.n112 iovss.n111 0.818682
R1911 iovss.n66 iovss.n64 0.818682
R1912 iovss.n117 iovss.n116 0.818682
R1913 iovss.n60 iovss.n59 0.818682
R1914 iovss.n127 iovss.n126 0.818682
R1915 iovss.n57 iovss.n55 0.818682
R1916 iovss.n132 iovss.n131 0.818682
R1917 iovss.n51 iovss.n50 0.818682
R1918 iovss.n142 iovss.n141 0.818682
R1919 iovss.n48 iovss.n46 0.818682
R1920 iovss.n147 iovss.n146 0.818682
R1921 iovss.n42 iovss.n41 0.818682
R1922 iovss.n157 iovss.n156 0.818682
R1923 iovss.n39 iovss.n37 0.818682
R1924 iovss.n162 iovss.n161 0.818682
R1925 iovss.n33 iovss.n32 0.818682
R1926 iovss.n172 iovss.n171 0.818682
R1927 iovss.n30 iovss.n28 0.818682
R1928 iovss.n177 iovss.n176 0.818682
R1929 iovss.n24 iovss.n23 0.818682
R1930 iovss.n187 iovss.n186 0.818682
R1931 iovss.n21 iovss.n19 0.818682
R1932 iovss.n192 iovss.n191 0.818682
R1933 iovss.n15 iovss.n14 0.818682
R1934 iovss.n202 iovss.n201 0.818682
R1935 iovss.n12 iovss.n10 0.818682
R1936 iovss.n207 iovss.n206 0.818682
R1937 iovss.n6 iovss.n5 0.818682
R1938 iovss.n217 iovss.n216 0.818682
R1939 iovss.n3 iovss.n2 0.818682
R1940 iovss.n85 iovss.n84 0.416993
R1941 iovss.n219 iovss.n218 0.416993
R1942 iovss.n90 iovss.n80 0.201704
R1943 iovss.n221 iovss.n220 0.2005
R1944 iovss.n215 iovss.n1 0.2005
R1945 iovss.n214 iovss.n213 0.2005
R1946 iovss.n11 iovss.n7 0.2005
R1947 iovss.n209 iovss.n208 0.2005
R1948 iovss.n200 iovss.n9 0.2005
R1949 iovss.n199 iovss.n198 0.2005
R1950 iovss.n20 iovss.n16 0.2005
R1951 iovss.n194 iovss.n193 0.2005
R1952 iovss.n185 iovss.n18 0.2005
R1953 iovss.n184 iovss.n183 0.2005
R1954 iovss.n29 iovss.n25 0.2005
R1955 iovss.n179 iovss.n178 0.2005
R1956 iovss.n170 iovss.n27 0.2005
R1957 iovss.n169 iovss.n168 0.2005
R1958 iovss.n38 iovss.n34 0.2005
R1959 iovss.n164 iovss.n163 0.2005
R1960 iovss.n155 iovss.n36 0.2005
R1961 iovss.n154 iovss.n153 0.2005
R1962 iovss.n47 iovss.n43 0.2005
R1963 iovss.n149 iovss.n148 0.2005
R1964 iovss.n140 iovss.n45 0.2005
R1965 iovss.n139 iovss.n138 0.2005
R1966 iovss.n56 iovss.n52 0.2005
R1967 iovss.n134 iovss.n133 0.2005
R1968 iovss.n125 iovss.n54 0.2005
R1969 iovss.n124 iovss.n123 0.2005
R1970 iovss.n65 iovss.n61 0.2005
R1971 iovss.n119 iovss.n118 0.2005
R1972 iovss.n110 iovss.n63 0.2005
R1973 iovss.n109 iovss.n108 0.2005
R1974 iovss.n74 iovss.n70 0.2005
R1975 iovss.n104 iovss.n103 0.2005
R1976 iovss.n95 iovss.n72 0.2005
R1977 iovss.n94 iovss.n93 0.2005
R1978 iovss.n82 iovss.n79 0.2005
R1979 iovss.n89 iovss.n88 0.2005
R1980 iovss.n222 iovss.n221 0.1105
R1981 iovss.n1 iovss.n0 0.1105
R1982 iovss.n213 iovss.n212 0.1105
R1983 iovss.n211 iovss.n7 0.1105
R1984 iovss.n210 iovss.n209 0.1105
R1985 iovss.n9 iovss.n8 0.1105
R1986 iovss.n198 iovss.n197 0.1105
R1987 iovss.n196 iovss.n16 0.1105
R1988 iovss.n195 iovss.n194 0.1105
R1989 iovss.n18 iovss.n17 0.1105
R1990 iovss.n183 iovss.n182 0.1105
R1991 iovss.n181 iovss.n25 0.1105
R1992 iovss.n180 iovss.n179 0.1105
R1993 iovss.n27 iovss.n26 0.1105
R1994 iovss.n168 iovss.n167 0.1105
R1995 iovss.n166 iovss.n34 0.1105
R1996 iovss.n165 iovss.n164 0.1105
R1997 iovss.n36 iovss.n35 0.1105
R1998 iovss.n153 iovss.n152 0.1105
R1999 iovss.n151 iovss.n43 0.1105
R2000 iovss.n150 iovss.n149 0.1105
R2001 iovss.n45 iovss.n44 0.1105
R2002 iovss.n138 iovss.n137 0.1105
R2003 iovss.n136 iovss.n52 0.1105
R2004 iovss.n135 iovss.n134 0.1105
R2005 iovss.n54 iovss.n53 0.1105
R2006 iovss.n123 iovss.n122 0.1105
R2007 iovss.n121 iovss.n61 0.1105
R2008 iovss.n120 iovss.n119 0.1105
R2009 iovss.n63 iovss.n62 0.1105
R2010 iovss.n108 iovss.n107 0.1105
R2011 iovss.n106 iovss.n70 0.1105
R2012 iovss.n105 iovss.n104 0.1105
R2013 iovss.n72 iovss.n71 0.1105
R2014 iovss.n93 iovss.n92 0.1105
R2015 iovss.n91 iovss.n79 0.1105
R2016 iovss.n91 iovss.n90 0.0568704
R2017 iovss.n85 iovss.n76 0.00740196
R2018 iovss.n98 iovss.n76 0.00740196
R2019 iovss.n99 iovss.n98 0.00740196
R2020 iovss.n100 iovss.n99 0.00740196
R2021 iovss.n100 iovss.n67 0.00740196
R2022 iovss.n113 iovss.n67 0.00740196
R2023 iovss.n114 iovss.n113 0.00740196
R2024 iovss.n115 iovss.n114 0.00740196
R2025 iovss.n115 iovss.n58 0.00740196
R2026 iovss.n128 iovss.n58 0.00740196
R2027 iovss.n129 iovss.n128 0.00740196
R2028 iovss.n130 iovss.n129 0.00740196
R2029 iovss.n130 iovss.n49 0.00740196
R2030 iovss.n143 iovss.n49 0.00740196
R2031 iovss.n144 iovss.n143 0.00740196
R2032 iovss.n145 iovss.n144 0.00740196
R2033 iovss.n145 iovss.n40 0.00740196
R2034 iovss.n158 iovss.n40 0.00740196
R2035 iovss.n159 iovss.n158 0.00740196
R2036 iovss.n160 iovss.n159 0.00740196
R2037 iovss.n160 iovss.n31 0.00740196
R2038 iovss.n173 iovss.n31 0.00740196
R2039 iovss.n174 iovss.n173 0.00740196
R2040 iovss.n175 iovss.n174 0.00740196
R2041 iovss.n175 iovss.n22 0.00740196
R2042 iovss.n188 iovss.n22 0.00740196
R2043 iovss.n189 iovss.n188 0.00740196
R2044 iovss.n190 iovss.n189 0.00740196
R2045 iovss.n190 iovss.n13 0.00740196
R2046 iovss.n203 iovss.n13 0.00740196
R2047 iovss.n204 iovss.n203 0.00740196
R2048 iovss.n205 iovss.n204 0.00740196
R2049 iovss.n205 iovss.n4 0.00740196
R2050 iovss.n218 iovss.n4 0.00740196
R2051 iovss.n86 iovss.n83 0.00740196
R2052 iovss.n86 iovss.n77 0.00740196
R2053 iovss.n97 iovss.n77 0.00740196
R2054 iovss.n97 iovss.n75 0.00740196
R2055 iovss.n101 iovss.n75 0.00740196
R2056 iovss.n101 iovss.n68 0.00740196
R2057 iovss.n112 iovss.n68 0.00740196
R2058 iovss.n112 iovss.n66 0.00740196
R2059 iovss.n116 iovss.n66 0.00740196
R2060 iovss.n116 iovss.n59 0.00740196
R2061 iovss.n127 iovss.n59 0.00740196
R2062 iovss.n127 iovss.n57 0.00740196
R2063 iovss.n131 iovss.n57 0.00740196
R2064 iovss.n131 iovss.n50 0.00740196
R2065 iovss.n142 iovss.n50 0.00740196
R2066 iovss.n142 iovss.n48 0.00740196
R2067 iovss.n146 iovss.n48 0.00740196
R2068 iovss.n146 iovss.n41 0.00740196
R2069 iovss.n157 iovss.n41 0.00740196
R2070 iovss.n157 iovss.n39 0.00740196
R2071 iovss.n161 iovss.n39 0.00740196
R2072 iovss.n161 iovss.n32 0.00740196
R2073 iovss.n172 iovss.n32 0.00740196
R2074 iovss.n172 iovss.n30 0.00740196
R2075 iovss.n176 iovss.n30 0.00740196
R2076 iovss.n176 iovss.n23 0.00740196
R2077 iovss.n187 iovss.n23 0.00740196
R2078 iovss.n187 iovss.n21 0.00740196
R2079 iovss.n191 iovss.n21 0.00740196
R2080 iovss.n191 iovss.n14 0.00740196
R2081 iovss.n202 iovss.n14 0.00740196
R2082 iovss.n202 iovss.n12 0.00740196
R2083 iovss.n206 iovss.n12 0.00740196
R2084 iovss.n206 iovss.n5 0.00740196
R2085 iovss.n217 iovss.n5 0.00740196
R2086 iovss.n217 iovss.n3 0.00740196
R2087 iovss.n219 iovss.n3 0.00442211
R2088 iovss.n84 iovss.n83 0.00442211
R2089 iovss.n81 iovss.n80 0.00395098
R2090 iovss.n88 iovss.n81 0.00395098
R2091 iovss.n88 iovss.n87 0.00395098
R2092 iovss.n87 iovss.n82 0.00395098
R2093 iovss.n82 iovss.n78 0.00395098
R2094 iovss.n94 iovss.n78 0.00395098
R2095 iovss.n96 iovss.n94 0.00395098
R2096 iovss.n96 iovss.n95 0.00395098
R2097 iovss.n95 iovss.n73 0.00395098
R2098 iovss.n103 iovss.n73 0.00395098
R2099 iovss.n103 iovss.n102 0.00395098
R2100 iovss.n102 iovss.n74 0.00395098
R2101 iovss.n74 iovss.n69 0.00395098
R2102 iovss.n109 iovss.n69 0.00395098
R2103 iovss.n111 iovss.n109 0.00395098
R2104 iovss.n111 iovss.n110 0.00395098
R2105 iovss.n110 iovss.n64 0.00395098
R2106 iovss.n118 iovss.n64 0.00395098
R2107 iovss.n118 iovss.n117 0.00395098
R2108 iovss.n117 iovss.n65 0.00395098
R2109 iovss.n65 iovss.n60 0.00395098
R2110 iovss.n124 iovss.n60 0.00395098
R2111 iovss.n126 iovss.n124 0.00395098
R2112 iovss.n126 iovss.n125 0.00395098
R2113 iovss.n125 iovss.n55 0.00395098
R2114 iovss.n133 iovss.n55 0.00395098
R2115 iovss.n133 iovss.n132 0.00395098
R2116 iovss.n132 iovss.n56 0.00395098
R2117 iovss.n56 iovss.n51 0.00395098
R2118 iovss.n139 iovss.n51 0.00395098
R2119 iovss.n141 iovss.n139 0.00395098
R2120 iovss.n141 iovss.n140 0.00395098
R2121 iovss.n140 iovss.n46 0.00395098
R2122 iovss.n148 iovss.n46 0.00395098
R2123 iovss.n148 iovss.n147 0.00395098
R2124 iovss.n147 iovss.n47 0.00395098
R2125 iovss.n47 iovss.n42 0.00395098
R2126 iovss.n154 iovss.n42 0.00395098
R2127 iovss.n156 iovss.n154 0.00395098
R2128 iovss.n156 iovss.n155 0.00395098
R2129 iovss.n155 iovss.n37 0.00395098
R2130 iovss.n163 iovss.n37 0.00395098
R2131 iovss.n163 iovss.n162 0.00395098
R2132 iovss.n162 iovss.n38 0.00395098
R2133 iovss.n38 iovss.n33 0.00395098
R2134 iovss.n169 iovss.n33 0.00395098
R2135 iovss.n171 iovss.n169 0.00395098
R2136 iovss.n171 iovss.n170 0.00395098
R2137 iovss.n170 iovss.n28 0.00395098
R2138 iovss.n178 iovss.n28 0.00395098
R2139 iovss.n178 iovss.n177 0.00395098
R2140 iovss.n177 iovss.n29 0.00395098
R2141 iovss.n29 iovss.n24 0.00395098
R2142 iovss.n184 iovss.n24 0.00395098
R2143 iovss.n186 iovss.n184 0.00395098
R2144 iovss.n186 iovss.n185 0.00395098
R2145 iovss.n185 iovss.n19 0.00395098
R2146 iovss.n193 iovss.n19 0.00395098
R2147 iovss.n193 iovss.n192 0.00395098
R2148 iovss.n192 iovss.n20 0.00395098
R2149 iovss.n20 iovss.n15 0.00395098
R2150 iovss.n199 iovss.n15 0.00395098
R2151 iovss.n201 iovss.n199 0.00395098
R2152 iovss.n201 iovss.n200 0.00395098
R2153 iovss.n200 iovss.n10 0.00395098
R2154 iovss.n208 iovss.n10 0.00395098
R2155 iovss.n208 iovss.n207 0.00395098
R2156 iovss.n207 iovss.n11 0.00395098
R2157 iovss.n11 iovss.n6 0.00395098
R2158 iovss.n214 iovss.n6 0.00395098
R2159 iovss.n216 iovss.n214 0.00395098
R2160 iovss.n216 iovss.n215 0.00395098
R2161 iovss.n215 iovss.n2 0.00395098
R2162 iovss.n220 iovss.n2 0.00395098
R2163 iovss.n221 iovss 0.00261765
R2164 iovss iovss.n222 0.00196667
R2165 iovss.n89 iovss.n79 0.00191176
R2166 iovss.n93 iovss.n79 0.00191176
R2167 iovss.n93 iovss.n72 0.00191176
R2168 iovss.n104 iovss.n72 0.00191176
R2169 iovss.n104 iovss.n70 0.00191176
R2170 iovss.n108 iovss.n70 0.00191176
R2171 iovss.n108 iovss.n63 0.00191176
R2172 iovss.n119 iovss.n63 0.00191176
R2173 iovss.n119 iovss.n61 0.00191176
R2174 iovss.n123 iovss.n61 0.00191176
R2175 iovss.n123 iovss.n54 0.00191176
R2176 iovss.n134 iovss.n54 0.00191176
R2177 iovss.n134 iovss.n52 0.00191176
R2178 iovss.n138 iovss.n52 0.00191176
R2179 iovss.n138 iovss.n45 0.00191176
R2180 iovss.n149 iovss.n45 0.00191176
R2181 iovss.n149 iovss.n43 0.00191176
R2182 iovss.n153 iovss.n43 0.00191176
R2183 iovss.n153 iovss.n36 0.00191176
R2184 iovss.n164 iovss.n36 0.00191176
R2185 iovss.n164 iovss.n34 0.00191176
R2186 iovss.n168 iovss.n34 0.00191176
R2187 iovss.n168 iovss.n27 0.00191176
R2188 iovss.n179 iovss.n27 0.00191176
R2189 iovss.n179 iovss.n25 0.00191176
R2190 iovss.n183 iovss.n25 0.00191176
R2191 iovss.n183 iovss.n18 0.00191176
R2192 iovss.n194 iovss.n18 0.00191176
R2193 iovss.n194 iovss.n16 0.00191176
R2194 iovss.n198 iovss.n16 0.00191176
R2195 iovss.n198 iovss.n9 0.00191176
R2196 iovss.n209 iovss.n9 0.00191176
R2197 iovss.n209 iovss.n7 0.00191176
R2198 iovss.n213 iovss.n7 0.00191176
R2199 iovss.n213 iovss.n1 0.00191176
R2200 iovss.n221 iovss.n1 0.00191176
R2201 iovss.n90 iovss.n89 0.0016983
R2202 iovss.n92 iovss.n91 0.00147778
R2203 iovss.n92 iovss.n71 0.00147778
R2204 iovss.n105 iovss.n71 0.00147778
R2205 iovss.n106 iovss.n105 0.00147778
R2206 iovss.n107 iovss.n106 0.00147778
R2207 iovss.n107 iovss.n62 0.00147778
R2208 iovss.n120 iovss.n62 0.00147778
R2209 iovss.n121 iovss.n120 0.00147778
R2210 iovss.n122 iovss.n121 0.00147778
R2211 iovss.n122 iovss.n53 0.00147778
R2212 iovss.n135 iovss.n53 0.00147778
R2213 iovss.n136 iovss.n135 0.00147778
R2214 iovss.n137 iovss.n136 0.00147778
R2215 iovss.n137 iovss.n44 0.00147778
R2216 iovss.n150 iovss.n44 0.00147778
R2217 iovss.n151 iovss.n150 0.00147778
R2218 iovss.n152 iovss.n151 0.00147778
R2219 iovss.n152 iovss.n35 0.00147778
R2220 iovss.n165 iovss.n35 0.00147778
R2221 iovss.n166 iovss.n165 0.00147778
R2222 iovss.n167 iovss.n166 0.00147778
R2223 iovss.n167 iovss.n26 0.00147778
R2224 iovss.n180 iovss.n26 0.00147778
R2225 iovss.n181 iovss.n180 0.00147778
R2226 iovss.n182 iovss.n181 0.00147778
R2227 iovss.n182 iovss.n17 0.00147778
R2228 iovss.n195 iovss.n17 0.00147778
R2229 iovss.n196 iovss.n195 0.00147778
R2230 iovss.n197 iovss.n196 0.00147778
R2231 iovss.n197 iovss.n8 0.00147778
R2232 iovss.n210 iovss.n8 0.00147778
R2233 iovss.n211 iovss.n210 0.00147778
R2234 iovss.n212 iovss.n211 0.00147778
R2235 iovss.n212 iovss.n0 0.00147778
R2236 iovss.n222 iovss.n0 0.00147778
R2237 c2p_en.n2 c2p_en.t0 15.0005
R2238 c2p_en.n1 c2p_en.t1 15.0005
R2239 c2p_en.n4 c2p_en.n1 9.74312
R2240 c2p_en.n3 c2p_en.n2 9.22574
R2241 c2p_en.n0 c2p_en 9.10188
R2242 c2p_en.n2 c2p_en 2.16907
R2243 c2p_en.n1 c2p_en 2.16907
R2244 c2p_en.n4 c2p_en.n0 1.63153
R2245 c2p_en.n0 c2p_en 0.99754
R2246 c2p_en c2p_en.n4 0.0885
R2247 c2p_en.n3 c2p_en 0.0308448
R2248 c2p_en.n4 c2p_en.n3 0.0141552
R2249 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t3 21.2194
R2250 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n0 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t2 15.755
R2251 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n1 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n0 12.6797
R2252 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n0 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq 1.8683
R2253 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n3 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t0 1.73646
R2254 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n3 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n2 1.57533
R2255 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n2 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t1 1.43953
R2256 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n2 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n1 0.782552
R2257 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n3 0.753577
R2258 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n1 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq 0.0764524
R2259 c2p.n2 c2p.t1 15.0005
R2260 c2p.n1 c2p.t0 15.0005
R2261 c2p.n4 c2p.n1 12.0592
R2262 c2p.n3 c2p.n2 11.3445
R2263 c2p.n0 c2p 9.10188
R2264 c2p.n2 c2p 2.16907
R2265 c2p.n1 c2p 2.16907
R2266 c2p.n4 c2p.n0 0.404086
R2267 c2p.n0 c2p 0.28562
R2268 c2p c2p.n4 0.0885
R2269 c2p.n3 c2p 0.0308448
R2270 c2p.n4 c2p.n3 0.0141552
R2271 vdd.n35 vdd.n34 23.1683
R2272 vdd.n26 vdd.t1 17.0005
R2273 vdd.n28 vdd.t3 17.0005
R2274 vdd.n30 vdd.t8 17.0005
R2275 vdd.n23 vdd.t7 17.0005
R2276 vdd.n26 vdd.t0 11.3504
R2277 vdd.n33 vdd.t4 11.3229
R2278 vdd.n21 vdd.n15 8.45671
R2279 vdd.n18 vdd.n15 8.45671
R2280 vdd.n29 vdd.n24 5.65625
R2281 vdd.n27 vdd.n24 5.65625
R2282 vdd.n32 vdd.n31 5.64342
R2283 vdd.n22 vdd.n15 5.58952
R2284 vdd.n14 vdd.n13 3.57695
R2285 vdd.n37 vdd.n36 3.44123
R2286 vdd.n25 vdd.n24 2.83433
R2287 vdd.n20 vdd.t9 2.67724
R2288 vdd.n17 vdd.t6 2.67724
R2289 vdd.n38 vdd.n13 2.5353
R2290 vdd.n19 vdd.n15 2.23769
R2291 vdd.n36 vdd.n35 1.91595
R2292 vdd.n17 vdd.n16 1.89106
R2293 vdd.n16 vdd.n13 1.79777
R2294 vdd.n100 vdd.n99 1.50539
R2295 vdd.n1 vdd.n0 1.5005
R2296 vdd.n95 vdd.n94 1.5005
R2297 vdd.n93 vdd.n92 1.5005
R2298 vdd.n5 vdd.n4 1.5005
R2299 vdd.n87 vdd.n86 1.5005
R2300 vdd.n85 vdd.n84 1.5005
R2301 vdd.n9 vdd.n8 1.5005
R2302 vdd.n79 vdd.n78 1.5005
R2303 vdd.n77 vdd.n76 1.5005
R2304 vdd.n39 vdd.n12 1.5005
R2305 vdd.n71 vdd.n70 1.5005
R2306 vdd.n69 vdd.n68 1.5005
R2307 vdd.n43 vdd.n42 1.5005
R2308 vdd.n63 vdd.n62 1.5005
R2309 vdd.n61 vdd.n60 1.5005
R2310 vdd.n47 vdd.n46 1.5005
R2311 vdd.n55 vdd.n54 1.5005
R2312 vdd.n53 vdd.n52 1.5005
R2313 vdd.n19 vdd 0.719163
R2314 vdd.n101 vdd 0.6957
R2315 vdd.n20 vdd.n19 0.675725
R2316 vdd.n35 vdd.n22 0.319001
R2317 vdd.n99 vdd.n98 0.314786
R2318 vdd.n97 vdd.n96 0.314786
R2319 vdd.n3 vdd.n2 0.314786
R2320 vdd.n91 vdd.n90 0.314786
R2321 vdd.n89 vdd.n88 0.314786
R2322 vdd.n7 vdd.n6 0.314786
R2323 vdd.n83 vdd.n82 0.314786
R2324 vdd.n81 vdd.n80 0.314786
R2325 vdd.n11 vdd.n10 0.314786
R2326 vdd.n75 vdd.n74 0.314786
R2327 vdd.n73 vdd.n72 0.314786
R2328 vdd.n41 vdd.n40 0.314786
R2329 vdd.n67 vdd.n66 0.314786
R2330 vdd.n65 vdd.n64 0.314786
R2331 vdd.n45 vdd.n44 0.314786
R2332 vdd.n59 vdd.n58 0.314786
R2333 vdd.n57 vdd.n56 0.314786
R2334 vdd.n49 vdd.n48 0.314786
R2335 vdd vdd.n18 0.296488
R2336 vdd vdd.n21 0.296488
R2337 vdd.n22 vdd 0.232915
R2338 vdd.n50 vdd 0.217715
R2339 vdd.n51 vdd.n50 0.146103
R2340 vdd.n18 vdd.n17 0.105298
R2341 vdd.n21 vdd.n20 0.105298
R2342 vdd.n77 vdd.n38 0.0983261
R2343 vdd.n31 vdd 0.0934694
R2344 vdd.n38 vdd.n37 0.0897467
R2345 vdd.n31 vdd.n23 0.0756715
R2346 vdd.n14 vdd.t5 0.0742737
R2347 vdd.n27 vdd 0.0540006
R2348 vdd.n29 vdd.n28 0.0475075
R2349 vdd.n33 vdd 0.0474603
R2350 vdd.n34 vdd.n33 0.0360492
R2351 vdd.n52 vdd.n51 0.0354467
R2352 vdd.n30 vdd.n29 0.0348561
R2353 vdd.n28 vdd.n27 0.0333284
R2354 vdd.n51 vdd.n48 0.0314255
R2355 vdd vdd.n26 0.0199792
R2356 vdd vdd.n30 0.0199792
R2357 vdd.n23 vdd 0.0199792
R2358 vdd.n34 vdd 0.0115764
R2359 vdd.n54 vdd.n53 0.00921287
R2360 vdd.n54 vdd.n46 0.00921287
R2361 vdd.n61 vdd.n46 0.00921287
R2362 vdd.n62 vdd.n61 0.00921287
R2363 vdd.n62 vdd.n42 0.00921287
R2364 vdd.n69 vdd.n42 0.00921287
R2365 vdd.n70 vdd.n69 0.00921287
R2366 vdd.n70 vdd.n12 0.00921287
R2367 vdd.n77 vdd.n12 0.00921287
R2368 vdd.n78 vdd.n77 0.00921287
R2369 vdd.n78 vdd.n8 0.00921287
R2370 vdd.n85 vdd.n8 0.00921287
R2371 vdd.n86 vdd.n85 0.00921287
R2372 vdd.n86 vdd.n4 0.00921287
R2373 vdd.n93 vdd.n4 0.00921287
R2374 vdd.n94 vdd.n93 0.00921287
R2375 vdd.n94 vdd.n0 0.00921287
R2376 vdd.n100 vdd.n0 0.00921287
R2377 vdd.n37 vdd 0.00903111
R2378 vdd.n52 vdd.n49 0.00538889
R2379 vdd.n55 vdd.n49 0.00538889
R2380 vdd.n56 vdd.n55 0.00538889
R2381 vdd.n56 vdd.n47 0.00538889
R2382 vdd.n59 vdd.n47 0.00538889
R2383 vdd.n60 vdd.n59 0.00538889
R2384 vdd.n60 vdd.n45 0.00538889
R2385 vdd.n63 vdd.n45 0.00538889
R2386 vdd.n64 vdd.n63 0.00538889
R2387 vdd.n64 vdd.n43 0.00538889
R2388 vdd.n67 vdd.n43 0.00538889
R2389 vdd.n68 vdd.n67 0.00538889
R2390 vdd.n68 vdd.n41 0.00538889
R2391 vdd.n71 vdd.n41 0.00538889
R2392 vdd.n72 vdd.n71 0.00538889
R2393 vdd.n72 vdd.n39 0.00538889
R2394 vdd.n75 vdd.n39 0.00538889
R2395 vdd.n76 vdd.n75 0.00538889
R2396 vdd.n76 vdd.n11 0.00538889
R2397 vdd.n79 vdd.n11 0.00538889
R2398 vdd.n80 vdd.n79 0.00538889
R2399 vdd.n80 vdd.n9 0.00538889
R2400 vdd.n83 vdd.n9 0.00538889
R2401 vdd.n84 vdd.n83 0.00538889
R2402 vdd.n84 vdd.n7 0.00538889
R2403 vdd.n87 vdd.n7 0.00538889
R2404 vdd.n88 vdd.n87 0.00538889
R2405 vdd.n88 vdd.n5 0.00538889
R2406 vdd.n91 vdd.n5 0.00538889
R2407 vdd.n92 vdd.n91 0.00538889
R2408 vdd.n92 vdd.n3 0.00538889
R2409 vdd.n95 vdd.n3 0.00538889
R2410 vdd.n96 vdd.n95 0.00538889
R2411 vdd.n96 vdd.n1 0.00538889
R2412 vdd.n99 vdd.n1 0.00538889
R2413 vdd.n53 vdd.n50 0.00485644
R2414 vdd.n101 vdd.n100 0.00485644
R2415 vdd vdd.n101 0.00485644
R2416 vdd.n98 vdd 0.0035
R2417 vdd.n57 vdd.n48 0.0025
R2418 vdd.n58 vdd.n57 0.0025
R2419 vdd.n58 vdd.n44 0.0025
R2420 vdd.n65 vdd.n44 0.0025
R2421 vdd.n66 vdd.n65 0.0025
R2422 vdd.n66 vdd.n40 0.0025
R2423 vdd.n73 vdd.n40 0.0025
R2424 vdd.n74 vdd.n73 0.0025
R2425 vdd.n74 vdd.n10 0.0025
R2426 vdd.n81 vdd.n10 0.0025
R2427 vdd.n82 vdd.n81 0.0025
R2428 vdd.n82 vdd.n6 0.0025
R2429 vdd.n89 vdd.n6 0.0025
R2430 vdd.n90 vdd.n89 0.0025
R2431 vdd.n90 vdd.n2 0.0025
R2432 vdd.n97 vdd.n2 0.0025
R2433 vdd.n98 vdd.n97 0.0025
R2434 vdd.n36 vdd.n15 0.00244471
R2435 vdd.n16 vdd.n15 0.00240956
R2436 vdd.n15 vdd.n14 0.00100215
R2437 vdd.n25 vdd.t2 0.001
R2438 vdd.t4 vdd.n32 0.001
R2439 vdd.t0 vdd.n25 0.001
R2440 vdd.n32 vdd.t2 0.001
C0 c2p sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq 0.56766f
C1 a_8358_31526# sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq 0.30586f
C2 pad iovdd 43.7879f
C3 vdd sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq 1.86758f
C4 a_7724_30170# sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq 0.1286f
C5 c2p_en sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq 1.6012f
C6 a_8358_30206# a_8426_30170# 0.37106f
C7 a_8358_30206# a_8358_31526# 0.15491f
C8 a_7724_30170# a_7656_30206# 0.37106f
C9 vdd a_7656_31526# 0.79589f
C10 a_7656_31526# sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq 0.99218f
C11 c2p c2p_en 0.53273f
C12 vdd sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq 1.00261f
C13 a_7656_30206# a_7656_31526# 0.15491f
C14 c2p sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq 0.43902f
C15 a_8426_30170# iovdd 0.84126f
C16 sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq 1.30685f
C17 sg13g2_DCNDiode_0.guard pad 7.46684f
C18 c2p_en sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq 1.59673f
C19 a_7724_30170# iovdd 0.84924f
C20 vdd c2p 1.52081f
C21 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq a_8426_30170# 0.1286f
C22 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq a_8358_31526# 0.99584f
C23 c2p sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq 0.65338f
C24 a_7656_30206# iovdd 0.30461f
C25 vdd c2p_en 1.46533f
C26 vdd sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq 2.09027f
C27 vdd a_8358_31526# 0.80342f
C28 a_8358_30206# iovdd 0.28407f
C29 pad iovss 0.12305p
C30 c2p_en iovss 2.18641f
C31 c2p iovss 2.43746f
C32 iovdd iovss 0.14269p
C33 vdd iovss 0.24688p
C34 a_8358_30206# iovss 0.23648f
C35 a_7656_30206# iovss 0.45339f
C36 a_8426_30170# iovss 1.28351f
C37 a_7724_30170# iovss 1.27718f
C38 a_8358_31526# iovss 1.34776f
C39 a_7656_31526# iovss 1.89714f
C40 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq iovss 3.01174f
C41 sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq iovss 2.75308f
C42 sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq iovss 1.32815f
C43 sg13g2_DCNDiode_0.guard iovss 53.69175f $ **FLOATING
C44 vdd.n38 iovss 0.41076f
C45 vdd.n48 iovss 0.31195f
C46 vdd.n50 iovss 0.27112f
C47 vdd.n51 iovss 0.24976f
C48 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t1 iovss 0.16985f
C49 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t3 iovss 0.12361f
C50 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t2 iovss 0.16083f
C51 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n0 iovss 0.78384f
C52 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t0 iovss 0.23765f
C53 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n3 iovss 0.5473f
C54 sg13g2_GateDecode_0.ngate.t1 iovss 0.13894f
C55 sg13g2_GateDecode_0.ngate.n0 iovss 0.1062f
C56 sg13g2_GateDecode_0.ngate.t0 iovss 0.27352f
C57 sg13g2_GateDecode_0.ngate.n1 iovss 0.22609f
C58 sg13g2_Clamp_N15N15D_0.gate iovss 5.27154f
C59 sg13g2_GateDecode_0.ngate.t3 iovss 0.58807f
C60 sg13g2_GateDecode_0.ngate.t15 iovss 0.57383f
C61 sg13g2_GateDecode_0.ngate.n2 iovss 0.31341f
C62 sg13g2_GateDecode_0.ngate.t11 iovss 0.57383f
C63 sg13g2_GateDecode_0.ngate.n3 iovss 0.1756f
C64 sg13g2_GateDecode_0.ngate.t5 iovss 0.57383f
C65 sg13g2_GateDecode_0.ngate.n4 iovss 0.1756f
C66 sg13g2_GateDecode_0.ngate.t9 iovss 0.57383f
C67 sg13g2_GateDecode_0.ngate.n5 iovss 0.1756f
C68 sg13g2_GateDecode_0.ngate.t8 iovss 0.57383f
C69 sg13g2_GateDecode_0.ngate.n6 iovss 0.1756f
C70 sg13g2_GateDecode_0.ngate.t16 iovss 0.57383f
C71 sg13g2_GateDecode_0.ngate.n7 iovss 0.1756f
C72 sg13g2_GateDecode_0.ngate.t6 iovss 0.57383f
C73 sg13g2_GateDecode_0.ngate.n8 iovss 0.1756f
C74 sg13g2_GateDecode_0.ngate.t17 iovss 0.57383f
C75 sg13g2_GateDecode_0.ngate.n9 iovss 0.1756f
C76 sg13g2_GateDecode_0.ngate.t14 iovss 0.57383f
C77 sg13g2_GateDecode_0.ngate.n10 iovss 0.1756f
C78 sg13g2_GateDecode_0.ngate.t4 iovss 0.57383f
C79 sg13g2_GateDecode_0.ngate.n11 iovss 0.1756f
C80 sg13g2_GateDecode_0.ngate.t13 iovss 0.57383f
C81 sg13g2_GateDecode_0.ngate.n12 iovss 0.1756f
C82 sg13g2_GateDecode_0.ngate.t7 iovss 0.57383f
C83 sg13g2_GateDecode_0.ngate.n13 iovss 0.1756f
C84 sg13g2_GateDecode_0.ngate.t2 iovss 0.57383f
C85 sg13g2_GateDecode_0.ngate.n14 iovss 0.1756f
C86 sg13g2_GateDecode_0.ngate.t10 iovss 0.57383f
C87 sg13g2_GateDecode_0.ngate.n15 iovss 0.36396f
C88 sg13g2_GateDecode_0.ngate.t12 iovss 0.11129f
C89 sg13g2_GateDecode_0.ngate.n16 iovss 0.2721f
C90 sg13g2_GateDecode_0.sg13g2_LevelUp_0.o iovss 3.83921f
C91 pad.t21 iovss 0.20342f
C92 pad.n0 iovss 0.19135f
C93 pad.n28 iovss 0.20626f
C94 pad.n29 iovss 0.20626f
C95 pad.n30 iovss 0.20626f
C96 pad.n31 iovss 0.20626f
C97 pad.n32 iovss 0.20626f
C98 pad.n33 iovss 0.20626f
C99 pad.n34 iovss 0.20626f
C100 pad.n35 iovss 0.20626f
C101 pad.n36 iovss 0.20626f
C102 pad.n37 iovss 0.20626f
C103 pad.n38 iovss 0.20626f
C104 pad.n39 iovss 0.20626f
C105 pad.n40 iovss 0.20626f
C106 pad.n41 iovss 0.20626f
C107 pad.n42 iovss 0.20626f
C108 pad.n43 iovss 0.20626f
C109 pad.n44 iovss 0.20626f
C110 pad.n45 iovss 0.20626f
C111 pad.n46 iovss 0.20626f
C112 pad.n47 iovss 0.20626f
C113 pad.n48 iovss 0.20626f
C114 pad.n49 iovss 0.20626f
C115 pad.n53 iovss 0.37242f
C116 pad.n55 iovss 0.10191f
C117 pad.n56 iovss 0.17404f
C118 pad.n62 iovss 0.37242f
C119 pad.n79 iovss 0.20626f
C120 pad.n80 iovss 0.20626f
C121 pad.n81 iovss 0.20626f
C122 pad.n82 iovss 0.20626f
C123 pad.n83 iovss 0.20626f
C124 pad.n84 iovss 0.20626f
C125 pad.n85 iovss 0.20626f
C126 pad.n86 iovss 0.20626f
C127 pad.n87 iovss 0.20626f
C128 pad.n88 iovss 0.20626f
C129 pad.n89 iovss 0.20626f
C130 pad.n90 iovss 0.20626f
C131 pad.n91 iovss 0.20626f
C132 pad.n92 iovss 0.20626f
C133 pad.n93 iovss 0.20626f
C134 pad.n94 iovss 0.20626f
C135 pad.n103 iovss 0.20626f
C136 pad.n104 iovss 0.20626f
C137 pad.n105 iovss 0.20626f
C138 pad.n106 iovss 0.20626f
C139 pad.n107 iovss 0.20626f
C140 pad.n108 iovss 0.20626f
C141 pad.n109 iovss 0.20626f
C142 pad.n118 iovss 0.20626f
C143 pad.n119 iovss 0.20626f
C144 pad.n120 iovss 0.20626f
C145 pad.n121 iovss 0.61199f
C146 pad.n122 iovss 0.20626f
C147 pad.n123 iovss 0.20626f
C148 pad.n124 iovss 0.20626f
C149 pad.n131 iovss 0.20709f
C150 pad.n132 iovss 0.20687f
C151 pad.n133 iovss 0.21243f
C152 pad.n134 iovss 0.20626f
C153 pad.n135 iovss 0.20626f
C154 pad.n136 iovss 0.20626f
C155 pad.n138 iovss 0.25885f
C156 pad.n139 iovss 0.31357f
C157 pad.n166 iovss 0.20626f
C158 pad.n167 iovss 0.20626f
C159 pad.n168 iovss 0.20626f
C160 pad.n169 iovss 0.20626f
C161 pad.n170 iovss 0.20626f
C162 pad.n171 iovss 0.20626f
C163 pad.n172 iovss 0.20626f
C164 pad.n173 iovss 0.20626f
C165 pad.n174 iovss 0.20626f
C166 pad.n203 iovss 0.20626f
C167 pad.n204 iovss 0.20626f
C168 pad.n205 iovss 0.20626f
C169 pad.n206 iovss 0.20626f
C170 pad.n207 iovss 0.20626f
C171 pad.n208 iovss 0.20626f
C172 pad.n209 iovss 0.20626f
C173 pad.n210 iovss 0.20626f
C174 pad.n211 iovss 0.20626f
C175 pad.n227 iovss 0.37572f
C176 pad.t24 iovss 1.21278f
C177 pad.t0 iovss 0.44346f
C178 pad.t2 iovss 0.31211f
C179 pad.n229 iovss 0.36724f
C180 pad.n230 iovss 0.12692f
C181 pad.n233 iovss 0.17404f
C182 pad.t9 iovss 0.44346f
C183 pad.t11 iovss 0.31211f
C184 pad.n238 iovss 0.36724f
C185 pad.n239 iovss 0.12692f
C186 pad.n241 iovss 0.14668f
C187 pad.t10 iovss 0.44346f
C188 pad.t1 iovss 0.31211f
C189 pad.n244 iovss 0.36724f
C190 pad.t12 iovss 0.44346f
C191 pad.t13 iovss 0.31211f
C192 pad.n246 iovss 0.36724f
C193 pad.n248 iovss 0.37242f
C194 pad.n249 iovss 0.12692f
C195 pad.t14 iovss 0.34274f
C196 pad.t15 iovss 0.21137f
C197 pad.n251 iovss 0.36723f
C198 pad.n252 iovss 0.13022f
C199 pad.n253 iovss 0.17404f
C200 pad.t4 iovss 0.44359f
C201 pad.t5 iovss 0.31211f
C202 pad.n256 iovss 0.36711f
C203 pad.n257 iovss 0.14668f
C204 pad.n261 iovss 0.10191f
C205 pad.n262 iovss 0.37242f
C206 pad.n263 iovss 0.10191f
C207 pad.n264 iovss 0.37242f
C208 pad.n265 iovss 0.12692f
C209 pad.n266 iovss 0.10191f
C210 pad.t7 iovss 0.44346f
C211 pad.t8 iovss 0.31211f
C212 pad.n269 iovss 0.36724f
C213 pad.t16 iovss 0.20342f
C214 pad.n270 iovss 0.19135f
C215 pad.n272 iovss 0.14668f
C216 pad.n274 iovss 0.37242f
C217 pad.n275 iovss 0.37242f
C218 pad.n276 iovss 0.12692f
C219 pad.t3 iovss 0.44346f
C220 pad.t6 iovss 0.31211f
C221 pad.n280 iovss 0.36724f
C222 pad.n282 iovss 0.37242f
C223 pad.n283 iovss 0.12692f
C224 pad.t26 iovss 1.21278f
C225 pad.n288 iovss 0.12692f
C226 pad.n290 iovss 0.37242f
C227 pad.t22 iovss 0.20342f
C228 pad.n295 iovss 0.19135f
C229 pad.t17 iovss 0.20342f
C230 pad.n316 iovss 0.19135f
C231 pad.n318 iovss 0.14668f
C232 pad.n319 iovss 0.37242f
C233 pad.n323 iovss 0.37242f
C234 pad.n324 iovss 0.37242f
C235 pad.t25 iovss 1.21278f
C236 pad.n329 iovss 0.37242f
C237 pad.t18 iovss 0.20342f
C238 pad.n330 iovss 0.19135f
C239 pad.n331 iovss 0.14668f
C240 pad.n332 iovss 0.37242f
C241 pad.n336 iovss 0.17404f
C242 pad.n337 iovss 0.37572f
C243 pad.n338 iovss 0.14998f
C244 pad.t23 iovss 0.13686f
C245 pad.n339 iovss 0.19136f
C246 pad.n357 iovss 0.20626f
C247 pad.n358 iovss 0.20626f
C248 pad.n359 iovss 0.20626f
C249 pad.n360 iovss 0.20626f
C250 pad.n361 iovss 0.20626f
C251 pad.n362 iovss 0.20626f
C252 pad.n363 iovss 0.20626f
C253 pad.n364 iovss 0.20626f
C254 pad.n365 iovss 0.20626f
C255 pad.n366 iovss 0.20626f
C256 pad.n367 iovss 0.20626f
C257 pad.n368 iovss 0.20626f
C258 pad.n369 iovss 0.20626f
C259 pad.n370 iovss 0.20626f
C260 pad.n371 iovss 0.20626f
C261 pad.n372 iovss 0.20626f
C262 pad.n373 iovss 0.20626f
C263 pad.n374 iovss 0.20626f
C264 pad.n375 iovss 0.20626f
C265 pad.n376 iovss 0.20626f
C266 pad.t20 iovss 0.20342f
C267 pad.n405 iovss 0.19135f
C268 pad.n406 iovss 0.14668f
C269 pad.t27 iovss 1.21278f
C270 pad.n411 iovss 0.14668f
C271 pad.t19 iovss 0.20342f
C272 pad.n412 iovss 0.19135f
C273 pad.n430 iovss 0.20626f
C274 pad.n431 iovss 0.20626f
C275 pad.n432 iovss 0.20626f
C276 pad.n433 iovss 0.20626f
C277 pad.n434 iovss 0.20626f
C278 pad.n435 iovss 0.20626f
C279 pad.n436 iovss 0.20626f
C280 pad.n437 iovss 0.20626f
C281 pad.n438 iovss 0.20626f
C282 pad.n439 iovss 0.20626f
C283 pad.n440 iovss 0.20626f
C284 pad.n441 iovss 0.20626f
C285 pad.n442 iovss 0.20626f
C286 pad.n443 iovss 0.20626f
C287 pad.n444 iovss 0.20626f
C288 pad.n445 iovss 0.20626f
C289 pad.n446 iovss 0.20626f
C290 pad.n447 iovss 0.20626f
C291 pad.n448 iovss 0.20626f
C292 pad.n449 iovss 0.20626f
C293 pad.n450 iovss 0.20626f
C294 pad.n451 iovss 0.20626f
C295 pad.n452 iovss 0.20626f
C296 pad.n453 iovss 0.20626f
C297 pad.n454 iovss 0.20626f
C298 pad.n455 iovss 0.20626f
C299 pad.n456 iovss 0.20626f
C300 pad.n457 iovss 0.20626f
C301 pad.n458 iovss 0.20626f
C302 pad.n459 iovss 0.31357f
C303 pad.n476 iovss 0.20626f
C304 pad.n485 iovss 0.25883f
C305 pad.n486 iovss 0.20709f
C306 pad.n487 iovss 0.20626f
C307 pad.n488 iovss 0.15469f
C308 pad.n489 iovss 0.20626f
C309 pad.n490 iovss 0.20626f
C310 pad.n491 iovss 0.20626f
C311 pad.n492 iovss 0.20626f
C312 pad.n493 iovss 0.20626f
C313 pad.n494 iovss 0.20626f
C314 pad.n495 iovss 0.20626f
C315 pad.n496 iovss 0.20626f
C316 pad.n497 iovss 0.20626f
C317 iovdd.t0 iovss 10.6688f
C318 iovdd.n75 iovss 0.50524f
C319 iovdd.n121 iovss 0.31308f
C320 iovdd.n122 iovss 0.41468f
C321 iovdd.n123 iovss 0.41468f
C322 iovdd.n124 iovss 0.41468f
C323 iovdd.n125 iovss 0.20734f
C324 iovdd.n126 iovss 0.20734f
C325 iovdd.n127 iovss 0.41468f
C326 iovdd.n128 iovss 0.36589f
C327 iovdd.n129 iovss 0.41468f
C328 iovdd.n130 iovss 0.20734f
C329 iovdd.n131 iovss 0.41468f
C330 iovdd.n132 iovss 0.28146f
C331 iovdd.n134 iovss 0.2058f
C332 iovdd.n135 iovss 0.41468f
C333 iovdd.n136 iovss 0.20734f
C334 iovdd.n137 iovss 0.20734f
C335 iovdd.n138 iovss 0.41468f
C336 iovdd.n139 iovss 0.36589f
C337 iovdd.n140 iovss 0.41468f
C338 iovdd.n141 iovss 0.20734f
C339 iovdd.n142 iovss 0.41468f
C340 iovdd.n143 iovss 0.31308f
C341 iovdd.n145 iovss 0.28976f
C342 iovdd.n146 iovss 0.41468f
C343 iovdd.n147 iovss 0.20734f
C344 iovdd.n148 iovss 0.20734f
C345 iovdd.n149 iovss 0.41468f
C346 iovdd.n150 iovss 0.36589f
C347 iovdd.n151 iovss 0.41468f
C348 iovdd.n152 iovss 0.20734f
C349 iovdd.n153 iovss 0.41468f
C350 iovdd.n154 iovss 0.41468f
C351 iovdd.n155 iovss 0.41468f
C352 iovdd.n156 iovss 0.20734f
C353 iovdd.n157 iovss 0.20734f
C354 iovdd.n158 iovss 0.41468f
C355 iovdd.n159 iovss 0.36589f
C356 iovdd.n160 iovss 0.41468f
C357 iovdd.n161 iovss 0.20734f
C358 iovdd.n162 iovss 0.41468f
C359 iovdd.n163 iovss 0.41468f
C360 iovdd.n164 iovss 0.41468f
C361 iovdd.n165 iovss 0.20734f
C362 iovdd.n166 iovss 0.20734f
C363 iovdd.n167 iovss 0.41468f
C364 iovdd.n168 iovss 0.36589f
C365 iovdd.n169 iovss 0.41468f
C366 iovdd.n170 iovss 0.20734f
C367 iovdd.n171 iovss 0.41468f
C368 iovdd.n172 iovss 0.41468f
C369 iovdd.n173 iovss 0.41468f
C370 iovdd.n174 iovss 0.20734f
C371 iovdd.n175 iovss 0.20734f
C372 iovdd.n176 iovss 0.41468f
C373 iovdd.n177 iovss 1.4382f
C374 iovdd.n178 iovss 0.41468f
C375 iovdd.n179 iovss 0.20734f
C376 iovdd.n180 iovss 0.41468f
C377 iovdd.n181 iovss 0.73153f
C378 iovdd.n182 iovss 0.20734f
C379 iovdd.n183 iovss 0.84973f
C380 iovdd.n184 iovss 0.41468f
C381 iovdd.n185 iovss 0.20734f
C382 iovdd.n186 iovss 0.20734f
C383 iovdd.n187 iovss 0.41468f
C384 iovdd.n188 iovss 0.64348f
C385 iovdd.n189 iovss 1.42908f
C386 iovdd.n190 iovss 0.41468f
C387 iovdd.n191 iovss 0.41468f
C388 iovdd.n192 iovss 0.20734f
C389 iovdd.n193 iovss 0.20734f
C390 iovdd.n194 iovss 0.20734f
C391 iovdd.n195 iovss 0.41468f
C392 iovdd.n196 iovss 0.36589f
C393 iovdd.n197 iovss 0.36589f
C394 iovdd.n198 iovss 0.36589f
C395 iovdd.n199 iovss 0.41468f
C396 iovdd.n200 iovss 0.20734f
C397 iovdd.n201 iovss 0.20734f
C398 iovdd.n202 iovss 0.41468f
C399 iovdd.n203 iovss 0.41468f
C400 iovdd.n204 iovss 0.41468f
C401 iovdd.n205 iovss 0.41468f
C402 iovdd.n206 iovss 0.41468f
C403 iovdd.n207 iovss 0.20734f
C404 iovdd.n208 iovss 0.20734f
C405 iovdd.n209 iovss 0.20734f
C406 iovdd.n210 iovss 0.41468f
C407 iovdd.n211 iovss 0.36589f
C408 iovdd.n212 iovss 0.36589f
C409 iovdd.n213 iovss 0.36589f
C410 iovdd.n214 iovss 0.41468f
C411 iovdd.n215 iovss 0.20734f
C412 iovdd.n216 iovss 0.20734f
C413 iovdd.n217 iovss 0.41468f
C414 iovdd.n218 iovss 0.41468f
C415 iovdd.n219 iovss 0.41468f
C416 iovdd.n220 iovss 0.41468f
C417 iovdd.n221 iovss 0.41468f
C418 iovdd.n222 iovss 0.20734f
C419 iovdd.n223 iovss 0.20734f
C420 iovdd.n224 iovss 0.20734f
C421 iovdd.n225 iovss 0.41468f
C422 iovdd.n226 iovss 0.36589f
C423 iovdd.n227 iovss 0.36589f
C424 iovdd.n228 iovss 0.36589f
C425 iovdd.n229 iovss 0.41468f
C426 iovdd.n230 iovss 0.20734f
C427 iovdd.n231 iovss 0.20734f
C428 iovdd.n232 iovss 0.41468f
C429 iovdd.n233 iovss 0.41468f
C430 iovdd.n234 iovss 0.22652f
C431 iovdd.n235 iovss 0.2058f
C432 iovdd.n237 iovss 0.17354f
C433 iovdd.n246 iovss 0.2058f
C434 iovdd.n247 iovss 0.31308f
C435 iovdd.n248 iovss 0.41468f
C436 iovdd.n249 iovss 0.20734f
C437 iovdd.n250 iovss 0.20734f
C438 iovdd.n251 iovss 0.20734f
C439 iovdd.n252 iovss 0.41468f
C440 iovdd.n253 iovss 0.36589f
C441 iovdd.n254 iovss 0.36589f
C442 iovdd.n255 iovss 0.36589f
C443 iovdd.n256 iovss 0.41468f
C444 iovdd.n257 iovss 0.20734f
C445 iovdd.n258 iovss 0.20734f
C446 iovdd.n259 iovss 0.41468f
C447 iovdd.n260 iovss 0.23066f
C448 iovdd.n261 iovss 0.2058f
C449 iovdd.n280 iovss 0.2058f
C450 iovdd.n281 iovss 0.23481f
C451 iovdd.n282 iovss 0.28561f
C452 iovdd.n283 iovss 0.41468f
C453 iovdd.n284 iovss 0.20734f
C454 iovdd.n285 iovss 0.20734f
C455 iovdd.n286 iovss 0.20734f
C456 iovdd.n287 iovss 0.41468f
C457 iovdd.n288 iovss 0.36589f
C458 iovdd.n289 iovss 0.36589f
C459 iovdd.n290 iovss 0.36589f
C460 iovdd.n291 iovss 0.41468f
C461 iovdd.n292 iovss 0.20734f
C462 iovdd.n293 iovss 0.20734f
C463 iovdd.n294 iovss 0.41468f
C464 iovdd.n295 iovss 0.31308f
C465 iovdd.n296 iovss 0.2058f
C466 iovdd.n307 iovss 0.2058f
C467 iovdd.n308 iovss 0.23896f
C468 iovdd.n309 iovss 0.41468f
C469 iovdd.n310 iovss 0.20734f
C470 iovdd.n311 iovss 0.20734f
C471 iovdd.n312 iovss 0.20734f
C472 iovdd.n313 iovss 0.41468f
C473 iovdd.n314 iovss 0.36589f
C474 iovdd.n315 iovss 0.36589f
C475 iovdd.n316 iovss 0.36589f
C476 iovdd.n317 iovss 0.36589f
C477 iovdd.n318 iovss 0.41468f
C478 iovdd.n319 iovss 0.20734f
C479 iovdd.n320 iovss 0.41468f
C480 iovdd.n321 iovss 0.41468f
C481 iovdd.n322 iovss 0.41468f
C482 iovdd.n323 iovss 0.20734f
C483 iovdd.n324 iovss 0.36589f
C484 iovdd.n325 iovss 0.36589f
C485 iovdd.n326 iovss 0.36589f
C486 iovdd.n327 iovss 0.41468f
C487 iovdd.n328 iovss 0.20734f
C488 iovdd.n329 iovss 0.41468f
C489 iovdd.n330 iovss 0.41468f
C490 iovdd.n331 iovss 0.41468f
C491 iovdd.n332 iovss 0.41468f
C492 iovdd.n333 iovss 0.20734f
C493 iovdd.n334 iovss 0.36589f
C494 iovdd.n335 iovss 0.36589f
C495 iovdd.n336 iovss 0.36589f
C496 iovdd.n337 iovss 0.41468f
C497 iovdd.n338 iovss 0.20734f
C498 iovdd.n339 iovss 0.41468f
C499 iovdd.n340 iovss 0.41468f
C500 iovdd.n341 iovss 0.41468f
C501 iovdd.n342 iovss 0.41468f
C502 iovdd.n343 iovss 0.20734f
C503 iovdd.n344 iovss 0.36589f
C504 iovdd.n345 iovss 0.36589f
C505 iovdd.n346 iovss 0.36589f
C506 iovdd.n347 iovss 0.41468f
C507 iovdd.n348 iovss 0.20734f
C508 iovdd.n349 iovss 0.41468f
C509 iovdd.n350 iovss 1.42908f
C510 iovdd.n351 iovss 0.64348f
C511 iovdd.n352 iovss 0.36589f
C512 iovdd.n353 iovss 0.45737f
C513 iovdd.n354 iovss 0.51835f
C514 iovdd.n355 iovss 0.72652f
C515 iovdd.n356 iovss 0.20734f
C516 iovdd.n357 iovss 0.41468f
C517 iovdd.n358 iovss 0.41468f
C518 iovdd.n359 iovss 0.20734f
C519 iovdd.n360 iovss 0.20734f
C520 iovdd.n361 iovss 0.41468f
C521 iovdd.n362 iovss 0.41468f
C522 iovdd.n363 iovss 0.20734f
C523 iovdd.n364 iovss 0.20734f
C524 iovdd.n365 iovss 0.41468f
C525 iovdd.n366 iovss 0.41468f
C526 iovdd.n367 iovss 0.20734f
C527 iovdd.n368 iovss 0.20734f
C528 iovdd.n369 iovss 0.41468f
C529 iovdd.n370 iovss 0.41468f
C530 iovdd.n371 iovss 0.20734f
C531 iovdd.n372 iovss 0.20734f
C532 iovdd.n373 iovss 0.41468f
C533 iovdd.n374 iovss 0.41468f
C534 iovdd.n375 iovss 0.20734f
C535 iovdd.n376 iovss 0.20734f
C536 iovdd.n377 iovss 0.41468f
C537 iovdd.n378 iovss 0.41468f
C538 iovdd.n379 iovss 0.20734f
C539 iovdd.n380 iovss 0.20734f
C540 iovdd.n381 iovss 0.41468f
C541 iovdd.n382 iovss 0.41468f
C542 iovdd.n383 iovss 0.20734f
C543 iovdd.n384 iovss 0.20734f
C544 iovdd.n385 iovss 0.41468f
C545 iovdd.n386 iovss 0.41468f
C546 iovdd.n387 iovss 0.20734f
C547 iovdd.n388 iovss 0.20734f
C548 iovdd.n389 iovss 0.41468f
C549 iovdd.n390 iovss 0.27732f
C550 iovdd.n391 iovss 0.2058f
C551 iovdd.n398 iovss 0.12423f
C552 iovdd.n400 iovss 0.19411f
C553 iovdd.n422 iovss 0.12707f
C554 iovdd.t31 iovss 3.20726f
C555 iovdd.n511 iovss 0.83155f
C556 sg13g2_GateDecode_0.pgate.t1 iovss 0.26498f
C557 sg13g2_GateDecode_0.pgate.n0 iovss 0.20255f
C558 sg13g2_GateDecode_0.pgate.t0 iovss 0.52165f
C559 sg13g2_GateDecode_0.pgate.n1 iovss 0.4312f
C560 sg13g2_GateDecode_0.pgate.t5 iovss 3.26396f
C561 sg13g2_GateDecode_0.pgate.t16 iovss 3.26396f
C562 sg13g2_GateDecode_0.pgate.t10 iovss 3.26396f
C563 sg13g2_GateDecode_0.pgate.t4 iovss 3.26396f
C564 sg13g2_GateDecode_0.pgate.t11 iovss 3.26396f
C565 sg13g2_GateDecode_0.pgate.t3 iovss 3.26396f
C566 sg13g2_GateDecode_0.pgate.t12 iovss 3.26396f
C567 sg13g2_GateDecode_0.pgate.t8 iovss 3.26396f
C568 sg13g2_GateDecode_0.pgate.t14 iovss 3.26396f
C569 sg13g2_GateDecode_0.pgate.t6 iovss 3.26396f
C570 sg13g2_GateDecode_0.pgate.t17 iovss 3.26396f
C571 sg13g2_GateDecode_0.pgate.t9 iovss 3.26396f
C572 sg13g2_GateDecode_0.pgate.t15 iovss 3.26396f
C573 sg13g2_GateDecode_0.pgate.t13 iovss 3.26396f
C574 sg13g2_GateDecode_0.pgate.t7 iovss 3.32677f
C575 sg13g2_GateDecode_0.pgate.n3 iovss 1.15191f
C576 sg13g2_GateDecode_0.pgate.n4 iovss 0.62981f
C577 sg13g2_GateDecode_0.pgate.n5 iovss 0.62981f
C578 sg13g2_GateDecode_0.pgate.n6 iovss 0.62981f
C579 sg13g2_GateDecode_0.pgate.n7 iovss 0.62981f
C580 sg13g2_GateDecode_0.pgate.n8 iovss 0.62981f
C581 sg13g2_GateDecode_0.pgate.n9 iovss 0.62981f
C582 sg13g2_GateDecode_0.pgate.n10 iovss 0.62981f
C583 sg13g2_GateDecode_0.pgate.n11 iovss 0.62981f
C584 sg13g2_GateDecode_0.pgate.n12 iovss 0.62981f
C585 sg13g2_GateDecode_0.pgate.n13 iovss 0.62981f
C586 sg13g2_GateDecode_0.pgate.n14 iovss 0.62981f
C587 sg13g2_GateDecode_0.pgate.n15 iovss 0.62981f
C588 sg13g2_GateDecode_0.pgate.n16 iovss 0.98205f
C589 sg13g2_GateDecode_0.pgate.t2 iovss 0.21106f
C590 sg13g2_GateDecode_0.pgate.n17 iovss 0.11367f
C591 sg13g2_GateDecode_0.pgate.n18 iovss 0.41088f
C592 sg13g2_GateDecode_0.pgate.n19 iovss 4.40844f
C593 sg13g2_GateDecode_0.sg13g2_LevelUp_1.o iovss 3.4918f
.ends

