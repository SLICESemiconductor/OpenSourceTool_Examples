* NGSPICE file created from sg13g2_IOPadIOVss_flat.ext - technology: ihp-sg13g2

.subckt sg13g2_IOPadIOVss_flat vdd iovss iovdd
X0 iovss iovdd dpantenna l=27.78u w=1.26u
X1 iovss iovdd dpantenna l=27.78u w=1.26u
X2 iovss iovss dantenna l=27.78u w=1.26u
X3 iovss iovss dantenna l=27.78u w=1.26u
C0 iovdd iovss 0.31051p
C1 vdd iovss 0.24621p
C2 sg13g2_DCNDiode_0.guard iovss 0.27183p $ **FLOATING
.ends

