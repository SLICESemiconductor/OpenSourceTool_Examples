* NGSPICE file created from sg13g2_IOPadVdd_flat.ext - technology: ihp-sg13g2

.subckt sg13g2_IOPadVdd_flat vdd vss iovdd iovss
X0 iovss sg13g2_RCClampInverter_0.out.t31 vdd.t117 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X1 vdd.t131 sg13g2_RCClampInverter_0.out.t32 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X2 vdd.t119 sg13g2_RCClampInverter_0.out.t33 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X3 vdd.t42 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t16 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X4 sg13g2_RCClampInverter_0.out.t5 sg13g2_RCClampInverter_0.in.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=1.71p ps=9.38u w=9u l=0.5u
X5 iovss sg13g2_RCClampInverter_0.out.t34 vdd.t89 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X6 iovss sg13g2_RCClampInverter_0.out.t35 vdd.t125 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X7 iovss sg13g2_RCClampInverter_0.out.t36 vdd.t88 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X8 vdd.t26 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t28 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X9 sg13g2_RCClampInverter_0.out.t4 sg13g2_RCClampInverter_0.in.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=1.71p ps=9.38u w=9u l=0.5u
X10 iovss sg13g2_RCClampInverter_0.out.t37 vdd.t86 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X11 iovss sg13g2_RCClampInverter_0.out.t38 vdd.t84 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X12 iovss sg13g2_RCClampInverter_0.out.t39 vdd.t138 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X13 vdd.t138 sg13g2_RCClampInverter_0.out.t40 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X14 iovss sg13g2_RCClampInverter_0.out.t41 vdd.t137 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X15 vdd.t113 sg13g2_RCClampInverter_0.out.t42 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X16 iovss sg13g2_RCClampInverter_0.out.t43 vdd.t80 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X17 vdd.t20 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t20 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X18 vdd.t28 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t19 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X19 iovss sg13g2_RCClampInverter_0.out.t44 vdd.t120 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X20 vdd.t111 sg13g2_RCClampInverter_0.out.t45 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X21 iovss sg13g2_RCClampInverter_0.out.t46 vdd.t77 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X22 iovss sg13g2_RCClampInverter_0.out.t47 vdd.t135 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X23 iovss sg13g2_RCClampInverter_0.out.t48 vdd.t74 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X24 vdd.t109 sg13g2_RCClampInverter_0.out.t49 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X25 sg13g2_RCClampInverter_0.out.t23 sg13g2_RCClampInverter_0.in.t1 vdd.t19 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X26 a_11365_11542# a_11695_7456# iovss rppd l=20u w=1u
X27 vdd.t24 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t29 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X28 iovss sg13g2_RCClampInverter_0.out.t50 vdd.t70 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X29 sg13g2_RCClampInverter_0.out.t15 sg13g2_RCClampInverter_0.in.t1 vdd.t2 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X30 a_8725_11542# a_9055_7456# iovss rppd l=20u w=1u
X31 vdd.t130 sg13g2_RCClampInverter_0.out.t51 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X32 vdd.t129 sg13g2_RCClampInverter_0.out.t52 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X33 iovss sg13g2_RCClampInverter_0.out.t53 vdd.t105 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X34 a_10045_11542# a_9715_7456# iovss rppd l=20u w=1u
X35 vdd.t104 sg13g2_RCClampInverter_0.out.t54 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X36 iovss sg13g2_RCClampInverter_0.out.t55 vdd.t133 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X37 iovss sg13g2_RCClampInverter_0.out.t56 vdd.t103 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X38 vdd.t101 sg13g2_RCClampInverter_0.out.t57 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X39 vdd.t51 sg13g2_RCClampInverter_0.out.t58 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X40 iovss sg13g2_RCClampInverter_0.out.t59 vdd.t65 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X41 vdd.t33 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t24 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X42 iovss sg13g2_RCClampInverter_0.out.t60 vdd.t63 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X43 sg13g2_RCClampInverter_0.out.t21 sg13g2_RCClampInverter_0.in.t1 vdd.t42 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X44 iovss sg13g2_RCClampInverter_0.in.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=2.24759n ps=2.5228m w=9u l=9.5u
X45 iovss sg13g2_RCClampInverter_0.out.t61 vdd.t60 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X46 iovss sg13g2_RCClampInverter_0.in.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X47 iovss sg13g2_RCClampInverter_0.out.t62 vdd.t96 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X48 a_4105_11542# a_4435_7456# iovss rppd l=20u w=1u
X49 a_7405_11542# a_7735_7456# iovss rppd l=20u w=1u
X50 vdd.t124 sg13g2_RCClampInverter_0.out.t63 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X51 vdd.t82 sg13g2_RCClampInverter_0.out.t64 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X52 iovss sg13g2_RCClampInverter_0.out.t31 vdd.t95 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X53 vdd.t137 sg13g2_RCClampInverter_0.out.t65 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X54 vdd.t136 sg13g2_RCClampInverter_0.out.t66 iovss iovss sg13_hv_nmos ad=3.256p pd=10.28u as=1.408p ps=5.04u w=4.4u l=0.6u
X55 iovss sg13g2_RCClampInverter_0.out.t34 vdd.t52 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X56 vdd.t123 sg13g2_RCClampInverter_0.out.t67 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X57 vdd.t122 sg13g2_RCClampInverter_0.out.t68 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X58 sg13g2_RCClampInverter_0.out.t30 sg13g2_RCClampInverter_0.in.t1 vdd.t8 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X59 sg13g2_RCClampInverter_0.out.t25 sg13g2_RCClampInverter_0.in.t1 vdd.t15 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X60 iovss sg13g2_RCClampInverter_0.out.t69 vdd.t92 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X61 iovss sg13g2_RCClampInverter_0.in.t2 sg13g2_RCClampInverter_0.out.t3 iovss sg13_hv_nmos ad=1.71p pd=9.38u as=1.71p ps=9.38u w=9u l=0.5u
X62 iovss sg13g2_RCClampInverter_0.out.t70 vdd.t64 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X63 iovss sg13g2_RCClampInverter_0.out.t71 vdd.t102 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X64 vdd.t135 sg13g2_RCClampInverter_0.out.t72 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X65 sg13g2_RCClampInverter_0.out.t12 sg13g2_RCClampInverter_0.in.t1 vdd.t14 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X66 iovss sg13g2_RCClampInverter_0.in.t2 sg13g2_RCClampInverter_0.out.t2 iovss sg13_hv_nmos ad=1.71p pd=9.38u as=1.71p ps=9.38u w=9u l=0.5u
X67 sg13g2_RCClampInverter_0.out.t16 sg13g2_RCClampInverter_0.in.t1 vdd.t13 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X68 iovss sg13g2_RCClampInverter_0.in.t2 sg13g2_RCClampInverter_0.out.t1 iovss sg13_hv_nmos ad=1.71p pd=9.38u as=1.71p ps=9.38u w=9u l=0.5u
X69 iovss sg13g2_RCClampInverter_0.in.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X70 iovss sg13g2_RCClampInverter_0.out.t73 vdd.t134 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X71 vdd.t118 sg13g2_RCClampInverter_0.out.t74 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X72 vdd.t116 sg13g2_RCClampInverter_0.out.t75 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X73 sg13g2_RCClampInverter_0.out.t14 sg13g2_RCClampInverter_0.in.t1 vdd.t12 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X74 iovss sg13g2_RCClampInverter_0.in.t2 sg13g2_RCClampInverter_0.out.t0 iovss sg13_hv_nmos ad=1.71p pd=9.38u as=1.71p ps=9.38u w=9u l=0.5u
X75 iovss sg13g2_RCClampInverter_0.in.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X76 vdd.t134 sg13g2_RCClampInverter_0.out.t76 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=2.068p ps=9.74u w=4.4u l=0.6u
X77 sg13g2_RCClampInverter_0.out.t7 sg13g2_RCClampInverter_0.in.t1 vdd.t11 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X78 iovss sg13g2_RCClampInverter_0.in.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X79 vdd.t115 sg13g2_RCClampInverter_0.out.t77 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X80 iovss sg13g2_RCClampInverter_0.out.t78 vdd.t83 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X81 a_4765_11542# a_5095_7456# iovss rppd l=20u w=1u
X82 a_8065_11542# a_8395_7456# iovss rppd l=20u w=1u
X83 vdd.t87 sg13g2_RCClampInverter_0.out.t45 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X84 vdd.t69 sg13g2_RCClampInverter_0.out.t79 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X85 vdd.t114 sg13g2_RCClampInverter_0.out.t80 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X86 iovss sg13g2_RCClampInverter_0.in.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X87 vdd.t66 sg13g2_RCClampInverter_0.out.t81 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X88 sg13g2_RCClampInverter_0.out.t11 sg13g2_RCClampInverter_0.in.t1 vdd.t22 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X89 vdd.t133 sg13g2_RCClampInverter_0.out.t82 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X90 sg13g2_RCClampInverter_0.out.t27 sg13g2_RCClampInverter_0.in.t1 vdd.t17 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X91 iovss sg13g2_RCClampInverter_0.out.t83 vdd.t132 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X92 sg13g2_RCClampInverter_0.out.t20 sg13g2_RCClampInverter_0.in.t1 vdd.t33 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X93 iovss sg13g2_RCClampInverter_0.in.t2 sg13g2_RCClampInverter_0.out.t5 iovss sg13_hv_nmos ad=1.71p pd=9.38u as=1.71p ps=9.38u w=9u l=0.5u
X94 vdd.t132 sg13g2_RCClampInverter_0.out.t84 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X95 iovss sg13g2_RCClampInverter_0.out.t85 vdd.t131 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X96 vdd.t112 sg13g2_RCClampInverter_0.out.t86 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X97 sg13g2_RCClampInverter_0.out.t9 sg13g2_RCClampInverter_0.in.t1 vdd.t16 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X98 sg13g2_RCClampInverter_0.out.t18 sg13g2_RCClampInverter_0.in.t1 vdd.t7 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X99 iovss sg13g2_RCClampInverter_0.in.t2 sg13g2_RCClampInverter_0.out.t4 iovss sg13_hv_nmos ad=1.71p pd=9.38u as=1.71p ps=9.38u w=9u l=0.5u
X100 vdd.t110 sg13g2_RCClampInverter_0.out.t52 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X101 vdd.t61 sg13g2_RCClampInverter_0.out.t87 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X102 vdd.t76 sg13g2_RCClampInverter_0.out.t54 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X103 a_10705_11542# a_11035_7456# iovss rppd l=20u w=1u
X104 vdd.t97 sg13g2_RCClampInverter_0.out.t88 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X105 sg13g2_RCClampInverter_0.out.t13 sg13g2_RCClampInverter_0.in.t1 vdd.t5 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X106 vdd.t108 sg13g2_RCClampInverter_0.out.t89 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X107 sg13g2_RCClampInverter_0.out.t26 sg13g2_RCClampInverter_0.in.t1 vdd.t1 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X108 vdd.t139 a_3775_7456# iovss rppd l=20u w=1u
X109 iovss sg13g2_RCClampInverter_0.out.t90 vdd.t85 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X110 sg13g2_RCClampInverter_0.out.t17 sg13g2_RCClampInverter_0.in.t1 vdd.t28 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X111 iovss sg13g2_RCClampInverter_0.out.t37 vdd.t130 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X112 iovss sg13g2_RCClampInverter_0.out.t91 vdd.t129 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X113 sg13g2_RCClampInverter_0.out.t10 sg13g2_RCClampInverter_0.in.t1 vdd.t3 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X114 iovss sg13g2_RCClampInverter_0.out.t92 vdd.t128 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X115 sg13g2_RCClampInverter_0.out.t24 sg13g2_RCClampInverter_0.in.t1 vdd.t26 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X116 vdd.t128 sg13g2_RCClampInverter_0.out.t93 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X117 iovss sg13g2_RCClampInverter_0.out.t94 vdd.t126 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X118 a_5425_11542# a_5095_7456# iovss rppd l=20u w=1u
X119 a_8725_11542# a_8395_7456# iovss rppd l=20u w=1u
X120 vdd.t127 sg13g2_RCClampInverter_0.out.t66 iovss iovss sg13_hv_nmos ad=3.256p pd=10.28u as=1.408p ps=5.04u w=4.4u l=0.6u
X121 vdd.t126 sg13g2_RCClampInverter_0.out.t95 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X122 vdd.t98 sg13g2_RCClampInverter_0.out.t96 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X123 vdd.t99 sg13g2_RCClampInverter_0.out.t67 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X124 vdd.t125 sg13g2_RCClampInverter_0.out.t97 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X125 iovss sg13g2_RCClampInverter_0.out.t44 vdd.t75 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X126 iovss sg13g2_RCClampInverter_0.out.t48 vdd.t124 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X127 iovss sg13g2_RCClampInverter_0.out.t98 vdd.t107 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X128 iovss sg13g2_RCClampInverter_0.out.t71 vdd.t72 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X129 vdd.t57 sg13g2_RCClampInverter_0.out.t33 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X130 sg13g2_RCClampInverter_0.out.t6 sg13g2_RCClampInverter_0.in.t1 vdd.t25 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=2.38p ps=14.68u w=7u l=0.5u
X131 iovss sg13g2_RCClampInverter_0.in.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X132 iovss sg13g2_RCClampInverter_0.in.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X133 iovss sg13g2_RCClampInverter_0.out.t36 vdd.t123 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X134 iovss sg13g2_RCClampInverter_0.out.t73 vdd.t121 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X135 vdd.t94 sg13g2_RCClampInverter_0.out.t74 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X136 iovss sg13g2_RCClampInverter_0.out.t99 vdd.t122 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X137 vdd.t121 sg13g2_RCClampInverter_0.out.t76 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=2.068p ps=9.74u w=4.4u l=0.6u
X138 vdd.t93 sg13g2_RCClampInverter_0.out.t77 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X139 vdd.t120 sg13g2_RCClampInverter_0.out.t79 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X140 a_6085_11542# a_5755_7456# iovss rppd l=20u w=1u
X141 a_9385_11542# a_9055_7456# iovss rppd l=20u w=1u
X142 iovss sg13g2_RCClampInverter_0.out.t41 vdd.t100 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X143 iovss sg13g2_RCClampInverter_0.out.t56 vdd.t119 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X144 iovss sg13g2_RCClampInverter_0.out.t43 vdd.t118 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X145 vdd.t117 sg13g2_RCClampInverter_0.out.t42 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X146 iovss sg13g2_RCClampInverter_0.out.t60 vdd.t116 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X147 a_10045_11542# a_10375_7456# iovss rppd l=20u w=1u
X148 sg13g2_RCClampInverter_0.out.t28 sg13g2_RCClampInverter_0.in.t1 vdd.t24 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X149 iovss sg13g2_RCClampInverter_0.out.t46 vdd.t115 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X150 iovss sg13g2_RCClampInverter_0.out.t100 vdd.t59 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X151 sg13g2_RCClampInverter_0.out.t8 sg13g2_RCClampInverter_0.in.t1 vdd.t10 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X152 iovss sg13g2_RCClampInverter_0.out.t101 vdd.t114 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X153 vdd.t22 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t10 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X154 sg13g2_RCClampInverter_0.out.t22 sg13g2_RCClampInverter_0.in.t1 vdd.t9 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X155 vdd.t68 sg13g2_RCClampInverter_0.out.t88 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X156 iovss sg13g2_RCClampInverter_0.out.t31 vdd.t113 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X157 sg13g2_RCClampInverter_0.in.t0 a_11695_7456# iovss rppd l=20u w=1u
X158 iovss sg13g2_RCClampInverter_0.out.t90 vdd.t53 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X159 iovss sg13g2_RCClampInverter_0.out.t34 vdd.t112 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X160 vdd.t79 sg13g2_RCClampInverter_0.out.t51 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X161 sg13g2_RCClampInverter_0.out.t19 sg13g2_RCClampInverter_0.in.t1 vdd.t20 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X162 a_4765_11542# a_4435_7456# iovss rppd l=20u w=1u
X163 iovss sg13g2_RCClampInverter_0.out.t53 vdd.t111 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X164 iovss sg13g2_RCClampInverter_0.out.t91 vdd.t110 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X165 iovss sg13g2_RCClampInverter_0.out.t102 vdd.t109 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X166 vdd.t19 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t22 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X167 iovss sg13g2_RCClampInverter_0.out.t92 vdd.t106 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X168 iovss sg13g2_RCClampInverter_0.out.t103 vdd.t108 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X169 vdd.t107 sg13g2_RCClampInverter_0.out.t58 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X170 sg13g2_RCClampInverter_0.out.t29 sg13g2_RCClampInverter_0.in.t1 vdd.t6 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X171 vdd.t106 sg13g2_RCClampInverter_0.out.t93 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X172 a_9385_11542# a_9715_7456# iovss rppd l=20u w=1u
X173 iovss sg13g2_RCClampInverter_0.in.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X174 a_6085_11542# a_6415_7456# iovss rppd l=20u w=1u
X175 vdd.t105 sg13g2_RCClampInverter_0.out.t45 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X176 iovss sg13g2_RCClampInverter_0.in.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X177 a_10705_11542# a_10375_7456# iovss rppd l=20u w=1u
X178 iovss sg13g2_RCClampInverter_0.out.t98 vdd.t81 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X179 iovss sg13g2_RCClampInverter_0.out.t62 vdd.t104 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X180 vdd.t103 sg13g2_RCClampInverter_0.out.t33 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X181 vdd.t102 sg13g2_RCClampInverter_0.out.t64 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X182 vdd.t67 sg13g2_RCClampInverter_0.out.t63 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X183 iovss sg13g2_RCClampInverter_0.out.t104 vdd.t101 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X184 vdd.t100 sg13g2_RCClampInverter_0.out.t65 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X185 iovss sg13g2_RCClampInverter_0.out.t36 vdd.t99 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X186 iovss sg13g2_RCClampInverter_0.out.t105 vdd.t98 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X187 vdd.t17 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t21 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X188 iovss sg13g2_RCClampInverter_0.out.t70 vdd.t97 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X189 vdd.t58 sg13g2_RCClampInverter_0.out.t52 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X190 vdd.t16 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t8 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X191 vdd.t96 sg13g2_RCClampInverter_0.out.t54 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X192 iovss sg13g2_RCClampInverter_0.out.t41 vdd.t71 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X193 a_6745_11542# a_7075_7456# iovss rppd l=20u w=1u
X194 vdd.t95 sg13g2_RCClampInverter_0.out.t42 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X195 iovss sg13g2_RCClampInverter_0.out.t43 vdd.t94 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X196 vdd.t56 sg13g2_RCClampInverter_0.out.t75 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X197 vdd.t15 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t30 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X198 a_11365_11542# a_11035_7456# iovss rppd l=20u w=1u
X199 iovss sg13g2_RCClampInverter_0.out.t46 vdd.t93 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X200 vdd.t92 sg13g2_RCClampInverter_0.out.t106 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X201 sg13g2_RCClampInverter_0.out.t3 sg13g2_RCClampInverter_0.in.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=1.71p ps=9.38u w=9u l=0.5u
X202 iovss sg13g2_RCClampInverter_0.in.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X203 vdd.t14 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t18 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X204 sg13g2_RCClampInverter_0.out.t2 sg13g2_RCClampInverter_0.in.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=1.71p ps=9.38u w=9u l=0.5u
X205 iovss sg13g2_RCClampInverter_0.in.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X206 vdd.t13 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t15 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X207 sg13g2_RCClampInverter_0.out.t1 sg13g2_RCClampInverter_0.in.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=3.06p ps=18.68u w=9u l=0.5u
X208 iovss sg13g2_RCClampInverter_0.out.t83 vdd.t91 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X209 sg13g2_RCClampInverter_0.out.t0 sg13g2_RCClampInverter_0.in.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=3.06p ps=18.68u w=9u l=0.5u
X210 vdd.t91 sg13g2_RCClampInverter_0.out.t84 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X211 vdd.t90 sg13g2_RCClampInverter_0.out.t66 iovss iovss sg13_hv_nmos ad=3.256p pd=10.28u as=1.408p ps=5.04u w=4.4u l=0.6u
X212 vdd.t12 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t13 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X213 vdd.t89 sg13g2_RCClampInverter_0.out.t86 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X214 vdd.t88 sg13g2_RCClampInverter_0.out.t67 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X215 vdd.t11 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t26 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X216 vdd.t10 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t7 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X217 iovss sg13g2_RCClampInverter_0.out.t53 vdd.t87 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X218 vdd.t86 sg13g2_RCClampInverter_0.out.t51 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X219 vdd.t85 sg13g2_RCClampInverter_0.out.t87 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X220 vdd.t84 sg13g2_RCClampInverter_0.out.t107 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X221 a_5425_11542# a_5755_7456# iovss rppd l=20u w=1u
X222 vdd.t83 sg13g2_RCClampInverter_0.out.t108 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X223 iovss sg13g2_RCClampInverter_0.out.t71 vdd.t82 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X224 vdd.t9 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t11 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X225 vdd.t81 sg13g2_RCClampInverter_0.out.t58 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X226 vdd.t8 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t27 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X227 iovss sg13g2_RCClampInverter_0.in.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X228 vdd.t80 sg13g2_RCClampInverter_0.out.t74 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X229 iovss sg13g2_RCClampInverter_0.out.t73 vdd.t78 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X230 iovss sg13g2_RCClampInverter_0.out.t37 vdd.t79 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X231 iovss sg13g2_RCClampInverter_0.in.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X232 a_4105_11542# a_3775_7456# iovss rppd l=20u w=1u
X233 a_7405_11542# a_7075_7456# iovss rppd l=20u w=1u
X234 vdd.t78 sg13g2_RCClampInverter_0.out.t76 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=2.068p ps=9.74u w=4.4u l=0.6u
X235 vdd.t7 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t9 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X236 vdd.t77 sg13g2_RCClampInverter_0.out.t77 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X237 iovss sg13g2_RCClampInverter_0.out.t62 vdd.t76 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X238 vdd.t75 sg13g2_RCClampInverter_0.out.t79 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X239 vdd.t6 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t14 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X240 vdd.t74 sg13g2_RCClampInverter_0.out.t63 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X241 vdd.t73 sg13g2_RCClampInverter_0.out.t109 iovss iovss sg13_hv_nmos ad=3.256p pd=10.28u as=1.408p ps=5.04u w=4.4u l=0.6u
X242 vdd.t5 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t23 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X243 vdd.t72 sg13g2_RCClampInverter_0.out.t64 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X244 vdd.t71 sg13g2_RCClampInverter_0.out.t65 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X245 vdd.t70 sg13g2_RCClampInverter_0.out.t110 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X246 vdd.t4 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t17 vdd.t0 sg13_hv_pmos ad=2.38p pd=14.68u as=1.33p ps=7.38u w=7u l=0.5u
X247 iovss sg13g2_RCClampInverter_0.out.t44 vdd.t69 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X248 iovss sg13g2_RCClampInverter_0.out.t70 vdd.t68 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X249 iovss sg13g2_RCClampInverter_0.out.t48 vdd.t67 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X250 iovss sg13g2_RCClampInverter_0.out.t111 vdd.t66 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X251 vdd.t3 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t12 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X252 vdd.t65 sg13g2_RCClampInverter_0.out.t112 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X253 vdd.t64 sg13g2_RCClampInverter_0.out.t88 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X254 a_8065_11542# a_7735_7456# iovss rppd l=20u w=1u
X255 iovss sg13g2_RCClampInverter_0.out.t113 vdd.t62 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X256 vdd.t63 sg13g2_RCClampInverter_0.out.t75 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X257 vdd.t62 sg13g2_RCClampInverter_0.out.t114 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=2.068p ps=9.74u w=4.4u l=0.6u
X258 iovss sg13g2_RCClampInverter_0.out.t90 vdd.t61 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X259 vdd.t60 sg13g2_RCClampInverter_0.out.t115 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X260 vdd.t59 sg13g2_RCClampInverter_0.out.t116 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X261 iovss sg13g2_RCClampInverter_0.out.t91 vdd.t58 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X262 iovss sg13g2_RCClampInverter_0.out.t117 dantenna l=0.48u w=0.48u
X263 iovss sg13g2_RCClampInverter_0.out.t56 vdd.t57 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X264 iovss sg13g2_RCClampInverter_0.out.t92 vdd.t55 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X265 vdd.t2 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t6 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X266 iovss sg13g2_RCClampInverter_0.out.t60 vdd.t56 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X267 iovss sg13g2_RCClampInverter_0.out.t83 vdd.t54 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X268 vdd.t55 sg13g2_RCClampInverter_0.out.t93 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X269 vdd.t1 sg13g2_RCClampInverter_0.in.t1 sg13g2_RCClampInverter_0.out.t25 vdd.t0 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X270 vdd.t54 sg13g2_RCClampInverter_0.out.t84 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X271 vdd.t53 sg13g2_RCClampInverter_0.out.t87 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X272 vdd.t52 sg13g2_RCClampInverter_0.out.t86 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X273 a_6745_11542# a_6415_7456# iovss rppd l=20u w=1u
X274 iovss sg13g2_RCClampInverter_0.out.t98 vdd.t51 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
R0 sg13g2_RCClampInverter_0.out.n85 sg13g2_RCClampInverter_0.out.t117 17.2912
R1 sg13g2_RCClampInverter_0.out.n2 sg13g2_RCClampInverter_0.out.n0 6.58671
R2 sg13g2_RCClampInverter_0.out.n82 sg13g2_RCClampInverter_0.out.n81 5.73421
R3 sg13g2_RCClampInverter_0.out.n80 sg13g2_RCClampInverter_0.out.n79 5.73421
R4 sg13g2_RCClampInverter_0.out.n78 sg13g2_RCClampInverter_0.out.n77 5.73421
R5 sg13g2_RCClampInverter_0.out.n76 sg13g2_RCClampInverter_0.out.n75 5.73421
R6 sg13g2_RCClampInverter_0.out.n74 sg13g2_RCClampInverter_0.out.n73 5.73421
R7 sg13g2_RCClampInverter_0.out.n72 sg13g2_RCClampInverter_0.out.n71 5.73421
R8 sg13g2_RCClampInverter_0.out.n70 sg13g2_RCClampInverter_0.out.n69 5.73421
R9 sg13g2_RCClampInverter_0.out.n68 sg13g2_RCClampInverter_0.out.n67 5.73421
R10 sg13g2_RCClampInverter_0.out.n66 sg13g2_RCClampInverter_0.out.n65 5.73421
R11 sg13g2_RCClampInverter_0.out.n64 sg13g2_RCClampInverter_0.out.n63 5.73421
R12 sg13g2_RCClampInverter_0.out.n62 sg13g2_RCClampInverter_0.out.n61 5.73421
R13 sg13g2_RCClampInverter_0.out.n60 sg13g2_RCClampInverter_0.out.n59 5.73421
R14 sg13g2_RCClampInverter_0.out.n58 sg13g2_RCClampInverter_0.out.n57 5.73421
R15 sg13g2_RCClampInverter_0.out.n56 sg13g2_RCClampInverter_0.out.n55 5.73421
R16 sg13g2_RCClampInverter_0.out.n54 sg13g2_RCClampInverter_0.out.n53 5.73421
R17 sg13g2_RCClampInverter_0.out.n52 sg13g2_RCClampInverter_0.out.n51 5.73421
R18 sg13g2_RCClampInverter_0.out.n50 sg13g2_RCClampInverter_0.out.n49 5.73421
R19 sg13g2_RCClampInverter_0.out.n48 sg13g2_RCClampInverter_0.out.n47 5.73421
R20 sg13g2_RCClampInverter_0.out.n46 sg13g2_RCClampInverter_0.out.n45 5.73421
R21 sg13g2_RCClampInverter_0.out.n44 sg13g2_RCClampInverter_0.out.n43 5.73421
R22 sg13g2_RCClampInverter_0.out.n42 sg13g2_RCClampInverter_0.out.n41 5.73421
R23 sg13g2_RCClampInverter_0.out.n40 sg13g2_RCClampInverter_0.out.n39 5.73421
R24 sg13g2_RCClampInverter_0.out.n38 sg13g2_RCClampInverter_0.out.n37 5.73421
R25 sg13g2_RCClampInverter_0.out.n36 sg13g2_RCClampInverter_0.out.n35 5.73421
R26 sg13g2_RCClampInverter_0.out.n34 sg13g2_RCClampInverter_0.out.n33 5.73421
R27 sg13g2_RCClampInverter_0.out.n32 sg13g2_RCClampInverter_0.out.n31 5.73421
R28 sg13g2_RCClampInverter_0.out.n30 sg13g2_RCClampInverter_0.out.n29 5.73421
R29 sg13g2_RCClampInverter_0.out.n28 sg13g2_RCClampInverter_0.out.n27 5.73421
R30 sg13g2_RCClampInverter_0.out.n26 sg13g2_RCClampInverter_0.out.n25 5.73421
R31 sg13g2_RCClampInverter_0.out.n24 sg13g2_RCClampInverter_0.out.n23 5.73421
R32 sg13g2_RCClampInverter_0.out.n22 sg13g2_RCClampInverter_0.out.n21 5.73421
R33 sg13g2_RCClampInverter_0.out.n20 sg13g2_RCClampInverter_0.out.n19 5.73421
R34 sg13g2_RCClampInverter_0.out.n18 sg13g2_RCClampInverter_0.out.n17 5.73421
R35 sg13g2_RCClampInverter_0.out.n16 sg13g2_RCClampInverter_0.out.n15 5.73421
R36 sg13g2_RCClampInverter_0.out.n14 sg13g2_RCClampInverter_0.out.n13 5.73421
R37 sg13g2_RCClampInverter_0.out.n12 sg13g2_RCClampInverter_0.out.n11 5.73421
R38 sg13g2_RCClampInverter_0.out.n10 sg13g2_RCClampInverter_0.out.n9 5.73421
R39 sg13g2_RCClampInverter_0.out.n8 sg13g2_RCClampInverter_0.out.n7 5.73421
R40 sg13g2_RCClampInverter_0.out.n6 sg13g2_RCClampInverter_0.out.n5 5.73421
R41 sg13g2_RCClampInverter_0.out.n4 sg13g2_RCClampInverter_0.out.n3 5.73421
R42 sg13g2_RCClampInverter_0.out.n2 sg13g2_RCClampInverter_0.out.n1 5.73421
R43 sg13g2_RCClampInverter_0.out.n84 sg13g2_RCClampInverter_0.out.n83 5.73421
R44 sg13g2_RCClampInverter_0.out sg13g2_RCClampInverter_0.out.n85 4.50322
R45 sg13g2_RCClampInverter_0.out.n85 sg13g2_RCClampInverter_0.out.n84 2.48679
R46 sg13g2_RCClampInverter_0.out.n86 sg13g2_RCClampInverter_0.out.t17 1.72119
R47 sg13g2_RCClampInverter_0.out.n108 sg13g2_RCClampInverter_0.out.t15 1.69835
R48 sg13g2_RCClampInverter_0.out.n107 sg13g2_RCClampInverter_0.out.t16 1.69835
R49 sg13g2_RCClampInverter_0.out.n106 sg13g2_RCClampInverter_0.out.t21 1.69835
R50 sg13g2_RCClampInverter_0.out.n105 sg13g2_RCClampInverter_0.out.t27 1.69835
R51 sg13g2_RCClampInverter_0.out.n104 sg13g2_RCClampInverter_0.out.t30 1.69835
R52 sg13g2_RCClampInverter_0.out.n103 sg13g2_RCClampInverter_0.out.t25 1.69835
R53 sg13g2_RCClampInverter_0.out.n102 sg13g2_RCClampInverter_0.out.t26 1.69835
R54 sg13g2_RCClampInverter_0.out.n101 sg13g2_RCClampInverter_0.out.t7 1.69835
R55 sg13g2_RCClampInverter_0.out.n100 sg13g2_RCClampInverter_0.out.t8 1.69835
R56 sg13g2_RCClampInverter_0.out.n99 sg13g2_RCClampInverter_0.out.t9 1.69835
R57 sg13g2_RCClampInverter_0.out.n98 sg13g2_RCClampInverter_0.out.t18 1.69835
R58 sg13g2_RCClampInverter_0.out.n97 sg13g2_RCClampInverter_0.out.t12 1.69835
R59 sg13g2_RCClampInverter_0.out.n96 sg13g2_RCClampInverter_0.out.t10 1.69835
R60 sg13g2_RCClampInverter_0.out.n95 sg13g2_RCClampInverter_0.out.t11 1.69835
R61 sg13g2_RCClampInverter_0.out.n94 sg13g2_RCClampInverter_0.out.t22 1.69835
R62 sg13g2_RCClampInverter_0.out.n93 sg13g2_RCClampInverter_0.out.t23 1.69835
R63 sg13g2_RCClampInverter_0.out.n92 sg13g2_RCClampInverter_0.out.t13 1.69835
R64 sg13g2_RCClampInverter_0.out.n91 sg13g2_RCClampInverter_0.out.t14 1.69835
R65 sg13g2_RCClampInverter_0.out.n90 sg13g2_RCClampInverter_0.out.t29 1.69835
R66 sg13g2_RCClampInverter_0.out.n89 sg13g2_RCClampInverter_0.out.t28 1.69835
R67 sg13g2_RCClampInverter_0.out.n88 sg13g2_RCClampInverter_0.out.t24 1.69835
R68 sg13g2_RCClampInverter_0.out.n87 sg13g2_RCClampInverter_0.out.t20 1.69835
R69 sg13g2_RCClampInverter_0.out.n86 sg13g2_RCClampInverter_0.out.t19 1.69835
R70 sg13g2_RCClampInverter_0.out.n109 sg13g2_RCClampInverter_0.out.t6 1.69585
R71 sg13g2_RCClampInverter_0.out.n111 sg13g2_RCClampInverter_0.out.t5 1.44241
R72 sg13g2_RCClampInverter_0.out.n110 sg13g2_RCClampInverter_0.out.t0 1.43866
R73 sg13g2_RCClampInverter_0.out.n110 sg13g2_RCClampInverter_0.out.t4 1.43866
R74 sg13g2_RCClampInverter_0.out.n110 sg13g2_RCClampInverter_0.out.t2 1.43866
R75 sg13g2_RCClampInverter_0.out.n111 sg13g2_RCClampInverter_0.out.t1 1.43866
R76 sg13g2_RCClampInverter_0.out.n111 sg13g2_RCClampInverter_0.out.t3 1.43866
R77 sg13g2_RCClampInverter_0.out.n4 sg13g2_RCClampInverter_0.out.n2 1.22425
R78 sg13g2_RCClampInverter_0.out.n8 sg13g2_RCClampInverter_0.out.n6 1.22425
R79 sg13g2_RCClampInverter_0.out.n12 sg13g2_RCClampInverter_0.out.n10 1.22425
R80 sg13g2_RCClampInverter_0.out.n16 sg13g2_RCClampInverter_0.out.n14 1.22425
R81 sg13g2_RCClampInverter_0.out.n20 sg13g2_RCClampInverter_0.out.n18 1.22425
R82 sg13g2_RCClampInverter_0.out.n24 sg13g2_RCClampInverter_0.out.n22 1.22425
R83 sg13g2_RCClampInverter_0.out.n28 sg13g2_RCClampInverter_0.out.n26 1.22425
R84 sg13g2_RCClampInverter_0.out.n32 sg13g2_RCClampInverter_0.out.n30 1.22425
R85 sg13g2_RCClampInverter_0.out.n36 sg13g2_RCClampInverter_0.out.n34 1.22425
R86 sg13g2_RCClampInverter_0.out.n40 sg13g2_RCClampInverter_0.out.n38 1.22425
R87 sg13g2_RCClampInverter_0.out.n44 sg13g2_RCClampInverter_0.out.n42 1.22425
R88 sg13g2_RCClampInverter_0.out.n48 sg13g2_RCClampInverter_0.out.n46 1.22425
R89 sg13g2_RCClampInverter_0.out.n52 sg13g2_RCClampInverter_0.out.n50 1.22425
R90 sg13g2_RCClampInverter_0.out.n56 sg13g2_RCClampInverter_0.out.n54 1.22425
R91 sg13g2_RCClampInverter_0.out.n60 sg13g2_RCClampInverter_0.out.n58 1.22425
R92 sg13g2_RCClampInverter_0.out.n64 sg13g2_RCClampInverter_0.out.n62 1.22425
R93 sg13g2_RCClampInverter_0.out.n68 sg13g2_RCClampInverter_0.out.n66 1.22425
R94 sg13g2_RCClampInverter_0.out.n72 sg13g2_RCClampInverter_0.out.n70 1.22425
R95 sg13g2_RCClampInverter_0.out.n76 sg13g2_RCClampInverter_0.out.n74 1.22425
R96 sg13g2_RCClampInverter_0.out.n80 sg13g2_RCClampInverter_0.out.n78 1.22425
R97 sg13g2_RCClampInverter_0.out.n84 sg13g2_RCClampInverter_0.out.n82 1.22425
R98 sg13g2_RCClampInverter_0.out.n6 sg13g2_RCClampInverter_0.out.n4 0.853
R99 sg13g2_RCClampInverter_0.out.n10 sg13g2_RCClampInverter_0.out.n8 0.853
R100 sg13g2_RCClampInverter_0.out.n14 sg13g2_RCClampInverter_0.out.n12 0.853
R101 sg13g2_RCClampInverter_0.out.n18 sg13g2_RCClampInverter_0.out.n16 0.853
R102 sg13g2_RCClampInverter_0.out.n22 sg13g2_RCClampInverter_0.out.n20 0.853
R103 sg13g2_RCClampInverter_0.out.n26 sg13g2_RCClampInverter_0.out.n24 0.853
R104 sg13g2_RCClampInverter_0.out.n30 sg13g2_RCClampInverter_0.out.n28 0.853
R105 sg13g2_RCClampInverter_0.out.n34 sg13g2_RCClampInverter_0.out.n32 0.853
R106 sg13g2_RCClampInverter_0.out.n38 sg13g2_RCClampInverter_0.out.n36 0.853
R107 sg13g2_RCClampInverter_0.out.n42 sg13g2_RCClampInverter_0.out.n40 0.853
R108 sg13g2_RCClampInverter_0.out.n46 sg13g2_RCClampInverter_0.out.n44 0.853
R109 sg13g2_RCClampInverter_0.out.n50 sg13g2_RCClampInverter_0.out.n48 0.853
R110 sg13g2_RCClampInverter_0.out.n54 sg13g2_RCClampInverter_0.out.n52 0.853
R111 sg13g2_RCClampInverter_0.out.n58 sg13g2_RCClampInverter_0.out.n56 0.853
R112 sg13g2_RCClampInverter_0.out.n62 sg13g2_RCClampInverter_0.out.n60 0.853
R113 sg13g2_RCClampInverter_0.out.n66 sg13g2_RCClampInverter_0.out.n64 0.853
R114 sg13g2_RCClampInverter_0.out.n70 sg13g2_RCClampInverter_0.out.n68 0.853
R115 sg13g2_RCClampInverter_0.out.n74 sg13g2_RCClampInverter_0.out.n72 0.853
R116 sg13g2_RCClampInverter_0.out.n78 sg13g2_RCClampInverter_0.out.n76 0.853
R117 sg13g2_RCClampInverter_0.out.n82 sg13g2_RCClampInverter_0.out.n80 0.853
R118 sg13g2_RCClampInverter_0.out.n110 sg13g2_RCClampInverter_0.out.n109 0.332192
R119 sg13g2_RCClampInverter_0.out.n111 sg13g2_RCClampInverter_0.out.n110 0.119159
R120 sg13g2_RCClampInverter_0.out sg13g2_RCClampInverter_0.out.n111 0.0570714
R121 sg13g2_RCClampInverter_0.out.n87 sg13g2_RCClampInverter_0.out.n86 0.0233437
R122 sg13g2_RCClampInverter_0.out.n88 sg13g2_RCClampInverter_0.out.n87 0.0233437
R123 sg13g2_RCClampInverter_0.out.n89 sg13g2_RCClampInverter_0.out.n88 0.0233437
R124 sg13g2_RCClampInverter_0.out.n90 sg13g2_RCClampInverter_0.out.n89 0.0233437
R125 sg13g2_RCClampInverter_0.out.n91 sg13g2_RCClampInverter_0.out.n90 0.0233437
R126 sg13g2_RCClampInverter_0.out.n92 sg13g2_RCClampInverter_0.out.n91 0.0233437
R127 sg13g2_RCClampInverter_0.out.n93 sg13g2_RCClampInverter_0.out.n92 0.0233437
R128 sg13g2_RCClampInverter_0.out.n94 sg13g2_RCClampInverter_0.out.n93 0.0233437
R129 sg13g2_RCClampInverter_0.out.n95 sg13g2_RCClampInverter_0.out.n94 0.0233437
R130 sg13g2_RCClampInverter_0.out.n96 sg13g2_RCClampInverter_0.out.n95 0.0233437
R131 sg13g2_RCClampInverter_0.out.n97 sg13g2_RCClampInverter_0.out.n96 0.0233437
R132 sg13g2_RCClampInverter_0.out.n98 sg13g2_RCClampInverter_0.out.n97 0.0233437
R133 sg13g2_RCClampInverter_0.out.n99 sg13g2_RCClampInverter_0.out.n98 0.0233437
R134 sg13g2_RCClampInverter_0.out.n100 sg13g2_RCClampInverter_0.out.n99 0.0233437
R135 sg13g2_RCClampInverter_0.out.n101 sg13g2_RCClampInverter_0.out.n100 0.0233437
R136 sg13g2_RCClampInverter_0.out.n102 sg13g2_RCClampInverter_0.out.n101 0.0233437
R137 sg13g2_RCClampInverter_0.out.n103 sg13g2_RCClampInverter_0.out.n102 0.0233437
R138 sg13g2_RCClampInverter_0.out.n104 sg13g2_RCClampInverter_0.out.n103 0.0233437
R139 sg13g2_RCClampInverter_0.out.n105 sg13g2_RCClampInverter_0.out.n104 0.0233437
R140 sg13g2_RCClampInverter_0.out.n106 sg13g2_RCClampInverter_0.out.n105 0.0233437
R141 sg13g2_RCClampInverter_0.out.n107 sg13g2_RCClampInverter_0.out.n106 0.0233437
R142 sg13g2_RCClampInverter_0.out.n108 sg13g2_RCClampInverter_0.out.n107 0.0233437
R143 sg13g2_RCClampInverter_0.out.n109 sg13g2_RCClampInverter_0.out.n108 0.0233437
R144 sg13g2_RCClampInverter_0.out.n83 sg13g2_RCClampInverter_0.out.t76 0.001
R145 sg13g2_RCClampInverter_0.out.n83 sg13g2_RCClampInverter_0.out.t114 0.001
R146 sg13g2_RCClampInverter_0.out.n0 sg13g2_RCClampInverter_0.out.t66 0.001
R147 sg13g2_RCClampInverter_0.out.n0 sg13g2_RCClampInverter_0.out.t109 0.001
R148 sg13g2_RCClampInverter_0.out.n1 sg13g2_RCClampInverter_0.out.t70 0.001
R149 sg13g2_RCClampInverter_0.out.n1 sg13g2_RCClampInverter_0.out.t85 0.001
R150 sg13g2_RCClampInverter_0.out.n3 sg13g2_RCClampInverter_0.out.t88 0.001
R151 sg13g2_RCClampInverter_0.out.n3 sg13g2_RCClampInverter_0.out.t32 0.001
R152 sg13g2_RCClampInverter_0.out.n5 sg13g2_RCClampInverter_0.out.t37 0.001
R153 sg13g2_RCClampInverter_0.out.n5 sg13g2_RCClampInverter_0.out.t99 0.001
R154 sg13g2_RCClampInverter_0.out.n7 sg13g2_RCClampInverter_0.out.t51 0.001
R155 sg13g2_RCClampInverter_0.out.n7 sg13g2_RCClampInverter_0.out.t68 0.001
R156 sg13g2_RCClampInverter_0.out.n9 sg13g2_RCClampInverter_0.out.t60 0.001
R157 sg13g2_RCClampInverter_0.out.n9 sg13g2_RCClampInverter_0.out.t103 0.001
R158 sg13g2_RCClampInverter_0.out.n11 sg13g2_RCClampInverter_0.out.t75 0.001
R159 sg13g2_RCClampInverter_0.out.n11 sg13g2_RCClampInverter_0.out.t89 0.001
R160 sg13g2_RCClampInverter_0.out.n13 sg13g2_RCClampInverter_0.out.t98 0.001
R161 sg13g2_RCClampInverter_0.out.n13 sg13g2_RCClampInverter_0.out.t47 0.001
R162 sg13g2_RCClampInverter_0.out.n15 sg13g2_RCClampInverter_0.out.t58 0.001
R163 sg13g2_RCClampInverter_0.out.n15 sg13g2_RCClampInverter_0.out.t72 0.001
R164 sg13g2_RCClampInverter_0.out.n17 sg13g2_RCClampInverter_0.out.t53 0.001
R165 sg13g2_RCClampInverter_0.out.n17 sg13g2_RCClampInverter_0.out.t69 0.001
R166 sg13g2_RCClampInverter_0.out.n19 sg13g2_RCClampInverter_0.out.t45 0.001
R167 sg13g2_RCClampInverter_0.out.n19 sg13g2_RCClampInverter_0.out.t106 0.001
R168 sg13g2_RCClampInverter_0.out.n21 sg13g2_RCClampInverter_0.out.t36 0.001
R169 sg13g2_RCClampInverter_0.out.n21 sg13g2_RCClampInverter_0.out.t50 0.001
R170 sg13g2_RCClampInverter_0.out.n23 sg13g2_RCClampInverter_0.out.t67 0.001
R171 sg13g2_RCClampInverter_0.out.n23 sg13g2_RCClampInverter_0.out.t110 0.001
R172 sg13g2_RCClampInverter_0.out.n25 sg13g2_RCClampInverter_0.out.t56 0.001
R173 sg13g2_RCClampInverter_0.out.n25 sg13g2_RCClampInverter_0.out.t102 0.001
R174 sg13g2_RCClampInverter_0.out.n27 sg13g2_RCClampInverter_0.out.t33 0.001
R175 sg13g2_RCClampInverter_0.out.n27 sg13g2_RCClampInverter_0.out.t49 0.001
R176 sg13g2_RCClampInverter_0.out.n29 sg13g2_RCClampInverter_0.out.t34 0.001
R177 sg13g2_RCClampInverter_0.out.n29 sg13g2_RCClampInverter_0.out.t105 0.001
R178 sg13g2_RCClampInverter_0.out.n31 sg13g2_RCClampInverter_0.out.t86 0.001
R179 sg13g2_RCClampInverter_0.out.n31 sg13g2_RCClampInverter_0.out.t96 0.001
R180 sg13g2_RCClampInverter_0.out.n33 sg13g2_RCClampInverter_0.out.t41 0.001
R181 sg13g2_RCClampInverter_0.out.n33 sg13g2_RCClampInverter_0.out.t55 0.001
R182 sg13g2_RCClampInverter_0.out.n35 sg13g2_RCClampInverter_0.out.t65 0.001
R183 sg13g2_RCClampInverter_0.out.n35 sg13g2_RCClampInverter_0.out.t82 0.001
R184 sg13g2_RCClampInverter_0.out.n37 sg13g2_RCClampInverter_0.out.t62 0.001
R185 sg13g2_RCClampInverter_0.out.n37 sg13g2_RCClampInverter_0.out.t78 0.001
R186 sg13g2_RCClampInverter_0.out.n39 sg13g2_RCClampInverter_0.out.t54 0.001
R187 sg13g2_RCClampInverter_0.out.n39 sg13g2_RCClampInverter_0.out.t108 0.001
R188 sg13g2_RCClampInverter_0.out.n41 sg13g2_RCClampInverter_0.out.t46 0.001
R189 sg13g2_RCClampInverter_0.out.n41 sg13g2_RCClampInverter_0.out.t61 0.001
R190 sg13g2_RCClampInverter_0.out.n43 sg13g2_RCClampInverter_0.out.t77 0.001
R191 sg13g2_RCClampInverter_0.out.n43 sg13g2_RCClampInverter_0.out.t115 0.001
R192 sg13g2_RCClampInverter_0.out.n45 sg13g2_RCClampInverter_0.out.t31 0.001
R193 sg13g2_RCClampInverter_0.out.n45 sg13g2_RCClampInverter_0.out.t104 0.001
R194 sg13g2_RCClampInverter_0.out.n47 sg13g2_RCClampInverter_0.out.t42 0.001
R195 sg13g2_RCClampInverter_0.out.n47 sg13g2_RCClampInverter_0.out.t57 0.001
R196 sg13g2_RCClampInverter_0.out.n49 sg13g2_RCClampInverter_0.out.t48 0.001
R197 sg13g2_RCClampInverter_0.out.n49 sg13g2_RCClampInverter_0.out.t101 0.001
R198 sg13g2_RCClampInverter_0.out.n51 sg13g2_RCClampInverter_0.out.t63 0.001
R199 sg13g2_RCClampInverter_0.out.n51 sg13g2_RCClampInverter_0.out.t80 0.001
R200 sg13g2_RCClampInverter_0.out.n53 sg13g2_RCClampInverter_0.out.t90 0.001
R201 sg13g2_RCClampInverter_0.out.n53 sg13g2_RCClampInverter_0.out.t35 0.001
R202 sg13g2_RCClampInverter_0.out.n55 sg13g2_RCClampInverter_0.out.t87 0.001
R203 sg13g2_RCClampInverter_0.out.n55 sg13g2_RCClampInverter_0.out.t97 0.001
R204 sg13g2_RCClampInverter_0.out.n57 sg13g2_RCClampInverter_0.out.t43 0.001
R205 sg13g2_RCClampInverter_0.out.n57 sg13g2_RCClampInverter_0.out.t59 0.001
R206 sg13g2_RCClampInverter_0.out.n59 sg13g2_RCClampInverter_0.out.t74 0.001
R207 sg13g2_RCClampInverter_0.out.n59 sg13g2_RCClampInverter_0.out.t112 0.001
R208 sg13g2_RCClampInverter_0.out.n61 sg13g2_RCClampInverter_0.out.t92 0.001
R209 sg13g2_RCClampInverter_0.out.n61 sg13g2_RCClampInverter_0.out.t39 0.001
R210 sg13g2_RCClampInverter_0.out.n63 sg13g2_RCClampInverter_0.out.t93 0.001
R211 sg13g2_RCClampInverter_0.out.n63 sg13g2_RCClampInverter_0.out.t40 0.001
R212 sg13g2_RCClampInverter_0.out.n65 sg13g2_RCClampInverter_0.out.t44 0.001
R213 sg13g2_RCClampInverter_0.out.n65 sg13g2_RCClampInverter_0.out.t100 0.001
R214 sg13g2_RCClampInverter_0.out.n67 sg13g2_RCClampInverter_0.out.t79 0.001
R215 sg13g2_RCClampInverter_0.out.n67 sg13g2_RCClampInverter_0.out.t116 0.001
R216 sg13g2_RCClampInverter_0.out.n69 sg13g2_RCClampInverter_0.out.t83 0.001
R217 sg13g2_RCClampInverter_0.out.n69 sg13g2_RCClampInverter_0.out.t94 0.001
R218 sg13g2_RCClampInverter_0.out.n71 sg13g2_RCClampInverter_0.out.t84 0.001
R219 sg13g2_RCClampInverter_0.out.n71 sg13g2_RCClampInverter_0.out.t95 0.001
R220 sg13g2_RCClampInverter_0.out.n73 sg13g2_RCClampInverter_0.out.t71 0.001
R221 sg13g2_RCClampInverter_0.out.n73 sg13g2_RCClampInverter_0.out.t111 0.001
R222 sg13g2_RCClampInverter_0.out.n75 sg13g2_RCClampInverter_0.out.t64 0.001
R223 sg13g2_RCClampInverter_0.out.n75 sg13g2_RCClampInverter_0.out.t81 0.001
R224 sg13g2_RCClampInverter_0.out.n77 sg13g2_RCClampInverter_0.out.t91 0.001
R225 sg13g2_RCClampInverter_0.out.n77 sg13g2_RCClampInverter_0.out.t38 0.001
R226 sg13g2_RCClampInverter_0.out.n79 sg13g2_RCClampInverter_0.out.t52 0.001
R227 sg13g2_RCClampInverter_0.out.n79 sg13g2_RCClampInverter_0.out.t107 0.001
R228 sg13g2_RCClampInverter_0.out.n81 sg13g2_RCClampInverter_0.out.t73 0.001
R229 sg13g2_RCClampInverter_0.out.n81 sg13g2_RCClampInverter_0.out.t113 0.001
R230 vdd.n778 vdd.n10 25.498
R231 vdd.n10 vdd.t139 4.97569
R232 vdd.n410 vdd.n408 4.5146
R233 vdd.n780 vdd.n779 4.5005
R234 vdd.n12 vdd.n8 4.5005
R235 vdd.n759 vdd.n758 4.5005
R236 vdd.n743 vdd.n17 4.5005
R237 vdd.n751 vdd.n750 4.5005
R238 vdd.n720 vdd.n19 4.5005
R239 vdd.n712 vdd.n711 4.5005
R240 vdd.n694 vdd.n31 4.5005
R241 vdd.n703 vdd.n702 4.5005
R242 vdd.n37 vdd.n33 4.5005
R243 vdd.n670 vdd.n669 4.5005
R244 vdd.n650 vdd.n45 4.5005
R245 vdd.n658 vdd.n657 4.5005
R246 vdd.n62 vdd.n55 4.5005
R247 vdd.n624 vdd.n623 4.5005
R248 vdd.n622 vdd.n71 4.5005
R249 vdd.n588 vdd.n70 4.5005
R250 vdd.n614 vdd.n613 4.5005
R251 vdd.n77 vdd.n73 4.5005
R252 vdd.n568 vdd.n567 4.5005
R253 vdd.n507 vdd.n85 4.5005
R254 vdd.n514 vdd.n87 4.5005
R255 vdd.n522 vdd.n521 4.5005
R256 vdd.n530 vdd.n366 4.5005
R257 vdd.n538 vdd.n537 4.5005
R258 vdd.n373 vdd.n365 4.5005
R259 vdd.n468 vdd.n364 4.5005
R260 vdd.n461 vdd.n363 4.5005
R261 vdd.n455 vdd.n362 4.5005
R262 vdd.n447 vdd.n361 4.5005
R263 vdd.n439 vdd.n360 4.5005
R264 vdd.n428 vdd.n359 4.5005
R265 vdd.n401 vdd.n358 4.5005
R266 vdd.n412 vdd.n411 4.5005
R267 vdd.n410 vdd.n409 4.5005
R268 vdd.n411 vdd.n357 4.5005
R269 vdd.n553 vdd.n358 4.5005
R270 vdd.n552 vdd.n359 4.5005
R271 vdd.n551 vdd.n360 4.5005
R272 vdd.n549 vdd.n361 4.5005
R273 vdd.n546 vdd.n362 4.5005
R274 vdd.n545 vdd.n363 4.5005
R275 vdd.n542 vdd.n364 4.5005
R276 vdd.n541 vdd.n365 4.5005
R277 vdd.n539 vdd.n538 4.5005
R278 vdd.n366 vdd.n89 4.5005
R279 vdd.n521 vdd.n86 4.5005
R280 vdd.n562 vdd.n87 4.5005
R281 vdd.n563 vdd.n85 4.5005
R282 vdd.n567 vdd.n566 4.5005
R283 vdd.n73 vdd.n72 4.5005
R284 vdd.n617 vdd.n614 4.5005
R285 vdd.n618 vdd.n70 4.5005
R286 vdd.n622 vdd.n621 4.5005
R287 vdd.n623 vdd.n54 4.5005
R288 vdd.n660 vdd.n55 4.5005
R289 vdd.n659 vdd.n658 4.5005
R290 vdd.n46 vdd.n45 4.5005
R291 vdd.n669 vdd.n668 4.5005
R292 vdd.n33 vdd.n32 4.5005
R293 vdd.n704 vdd.n703 4.5005
R294 vdd.n707 vdd.n31 4.5005
R295 vdd.n711 vdd.n710 4.5005
R296 vdd.n19 vdd.n18 4.5005
R297 vdd.n752 vdd.n751 4.5005
R298 vdd.n755 vdd.n17 4.5005
R299 vdd.n758 vdd.n757 4.5005
R300 vdd.n8 vdd.n7 4.5005
R301 vdd.n781 vdd.n780 4.5005
R302 vdd.n266 vdd.n216 3.31474
R303 vdd.n266 vdd.n220 3.31474
R304 vdd.n266 vdd.n226 3.31474
R305 vdd.n266 vdd.n230 3.31474
R306 vdd.n266 vdd.n236 3.31474
R307 vdd.n266 vdd.n240 3.31474
R308 vdd.n266 vdd.n244 3.31474
R309 vdd.n266 vdd.n250 3.31474
R310 vdd.n266 vdd.n254 3.31474
R311 vdd.n266 vdd.n260 3.31474
R312 vdd.n266 vdd.n265 3.31474
R313 vdd.n266 vdd.n218 3.31457
R314 vdd.n266 vdd.n222 3.31457
R315 vdd.n266 vdd.n228 3.31457
R316 vdd.n266 vdd.n232 3.31457
R317 vdd.n266 vdd.n238 3.31457
R318 vdd.n266 vdd.n242 3.31457
R319 vdd.n266 vdd.n248 3.31457
R320 vdd.n266 vdd.n252 3.31457
R321 vdd.n266 vdd.n256 3.31457
R322 vdd.n266 vdd.n262 3.31457
R323 vdd.n257 vdd.t26 3.28171
R324 vdd.n223 vdd.t17 3.28171
R325 vdd.n263 vdd.t4 3.28171
R326 vdd.n264 vdd.t28 3.28171
R327 vdd.n261 vdd.t20 3.28171
R328 vdd.n259 vdd.t33 3.28171
R329 vdd.n255 vdd.t24 3.28171
R330 vdd.n253 vdd.t6 3.28171
R331 vdd.n251 vdd.t12 3.28171
R332 vdd.n249 vdd.t5 3.28171
R333 vdd.n247 vdd.t19 3.28171
R334 vdd.n245 vdd.t9 3.28171
R335 vdd.n243 vdd.t22 3.28171
R336 vdd.n241 vdd.t3 3.28171
R337 vdd.n239 vdd.t14 3.28171
R338 vdd.n237 vdd.t7 3.28171
R339 vdd.n235 vdd.t16 3.28171
R340 vdd.n233 vdd.t10 3.28171
R341 vdd.n231 vdd.t11 3.28171
R342 vdd.n229 vdd.t1 3.28171
R343 vdd.n227 vdd.t15 3.28171
R344 vdd.n225 vdd.t8 3.28171
R345 vdd.n221 vdd.t42 3.28171
R346 vdd.n219 vdd.t13 3.28171
R347 vdd.n217 vdd.t2 3.28171
R348 vdd.n215 vdd.t25 3.28171
R349 vdd.n266 vdd.n246 2.73027
R350 vdd.n266 vdd.n224 2.73011
R351 vdd.n266 vdd.n234 2.73011
R352 vdd.n266 vdd.n258 2.73011
R353 vdd.n397 vdd.t68 2.48354
R354 vdd.n433 vdd.t86 2.48354
R355 vdd.n388 vdd.t63 2.48354
R356 vdd.n381 vdd.t81 2.48354
R357 vdd.n376 vdd.t87 2.48354
R358 vdd.n369 vdd.t99 2.48354
R359 vdd.n487 vdd.t103 2.48354
R360 vdd.n494 vdd.t52 2.48354
R361 vdd.n500 vdd.t71 2.48354
R362 vdd.n78 vdd.t76 2.48354
R363 vdd.n584 vdd.t93 2.48354
R364 vdd.n591 vdd.t95 2.48354
R365 vdd.n65 vdd.t74 2.48354
R366 vdd.n58 vdd.t53 2.48354
R367 vdd.n643 vdd.t94 2.48354
R368 vdd.n38 vdd.t106 2.48354
R369 vdd.n686 vdd.t120 2.48354
R370 vdd.n26 vdd.t54 2.48354
R371 vdd.n724 vdd.t72 2.48354
R372 vdd.n736 vdd.t110 2.48354
R373 vdd.n763 vdd.t121 2.48354
R374 vdd.n404 vdd.t127 2.48325
R375 vdd.n409 vdd.n90 2.20698
R376 vdd.n782 vdd.n781 2.2005
R377 vdd.n7 vdd.n2 2.2005
R378 vdd.n757 vdd.n756 2.2005
R379 vdd.n755 vdd.n754 2.2005
R380 vdd.n753 vdd.n752 2.2005
R381 vdd.n708 vdd.n18 2.2005
R382 vdd.n710 vdd.n709 2.2005
R383 vdd.n707 vdd.n706 2.2005
R384 vdd.n705 vdd.n704 2.2005
R385 vdd.n666 vdd.n32 2.2005
R386 vdd.n668 vdd.n667 2.2005
R387 vdd.n665 vdd.n46 2.2005
R388 vdd.n659 vdd.n47 2.2005
R389 vdd.n661 vdd.n660 2.2005
R390 vdd.n54 vdd.n53 2.2005
R391 vdd.n621 vdd.n620 2.2005
R392 vdd.n619 vdd.n618 2.2005
R393 vdd.n617 vdd.n616 2.2005
R394 vdd.n615 vdd.n72 2.2005
R395 vdd.n566 vdd.n565 2.2005
R396 vdd.n564 vdd.n563 2.2005
R397 vdd.n562 vdd.n561 2.2005
R398 vdd.n560 vdd.n86 2.2005
R399 vdd.n559 vdd.n89 2.2005
R400 vdd.n539 vdd.n88 2.2005
R401 vdd.n541 vdd.n540 2.2005
R402 vdd.n543 vdd.n542 2.2005
R403 vdd.n545 vdd.n544 2.2005
R404 vdd.n547 vdd.n546 2.2005
R405 vdd.n549 vdd.n548 2.2005
R406 vdd.n551 vdd.n550 2.2005
R407 vdd.n552 vdd.n355 2.2005
R408 vdd.n554 vdd.n553 2.2005
R409 vdd.n357 vdd.n356 2.2005
R410 vdd.n397 vdd.t97 1.78531
R411 vdd.n398 vdd.t64 1.78531
R412 vdd.n399 vdd.t131 1.78531
R413 vdd.n433 vdd.t79 1.78531
R414 vdd.n434 vdd.t130 1.78531
R415 vdd.n435 vdd.t122 1.78531
R416 vdd.n388 vdd.t56 1.78531
R417 vdd.n389 vdd.t116 1.78531
R418 vdd.n390 vdd.t108 1.78531
R419 vdd.n381 vdd.t107 1.78531
R420 vdd.n382 vdd.t51 1.78531
R421 vdd.n383 vdd.t135 1.78531
R422 vdd.n376 vdd.t111 1.78531
R423 vdd.n377 vdd.t105 1.78531
R424 vdd.n378 vdd.t92 1.78531
R425 vdd.n369 vdd.t123 1.78531
R426 vdd.n370 vdd.t88 1.78531
R427 vdd.n371 vdd.t70 1.78531
R428 vdd.n487 vdd.t57 1.78531
R429 vdd.n488 vdd.t119 1.78531
R430 vdd.n489 vdd.t109 1.78531
R431 vdd.n494 vdd.t89 1.78531
R432 vdd.n495 vdd.t112 1.78531
R433 vdd.n496 vdd.t98 1.78531
R434 vdd.n500 vdd.t100 1.78531
R435 vdd.n501 vdd.t137 1.78531
R436 vdd.n502 vdd.t133 1.78531
R437 vdd.n78 vdd.t104 1.78531
R438 vdd.n79 vdd.t96 1.78531
R439 vdd.n80 vdd.t83 1.78531
R440 vdd.n584 vdd.t115 1.78531
R441 vdd.n585 vdd.t77 1.78531
R442 vdd.n586 vdd.t60 1.78531
R443 vdd.n591 vdd.t117 1.78531
R444 vdd.n592 vdd.t113 1.78531
R445 vdd.n593 vdd.t101 1.78531
R446 vdd.n65 vdd.t67 1.78531
R447 vdd.n66 vdd.t124 1.78531
R448 vdd.n67 vdd.t114 1.78531
R449 vdd.n58 vdd.t85 1.78531
R450 vdd.n59 vdd.t61 1.78531
R451 vdd.n60 vdd.t125 1.78531
R452 vdd.n643 vdd.t118 1.78531
R453 vdd.n644 vdd.t80 1.78531
R454 vdd.n645 vdd.t65 1.78531
R455 vdd.n38 vdd.t128 1.78531
R456 vdd.n39 vdd.t55 1.78531
R457 vdd.n40 vdd.t138 1.78531
R458 vdd.n686 vdd.t69 1.78531
R459 vdd.n687 vdd.t75 1.78531
R460 vdd.n688 vdd.t59 1.78531
R461 vdd.n26 vdd.t91 1.78531
R462 vdd.n27 vdd.t132 1.78531
R463 vdd.n28 vdd.t126 1.78531
R464 vdd.n724 vdd.t102 1.78531
R465 vdd.n725 vdd.t82 1.78531
R466 vdd.n726 vdd.t66 1.78531
R467 vdd.n736 vdd.t129 1.78531
R468 vdd.n737 vdd.t58 1.78531
R469 vdd.n738 vdd.t84 1.78531
R470 vdd.n763 vdd.t134 1.78531
R471 vdd.n764 vdd.t78 1.78531
R472 vdd.n765 vdd.t62 1.78531
R473 vdd.n404 vdd.t136 1.78502
R474 vdd.n405 vdd.t90 1.78502
R475 vdd.n406 vdd.t73 1.78502
R476 vdd.n290 vdd.n289 1.5005
R477 vdd.n287 vdd.n286 1.5005
R478 vdd.n294 vdd.n285 1.5005
R479 vdd.n297 vdd.n296 1.5005
R480 vdd.n299 vdd.n298 1.5005
R481 vdd.n302 vdd.n301 1.5005
R482 vdd.n304 vdd.n303 1.5005
R483 vdd.n284 vdd.n210 1.5005
R484 vdd.n283 vdd.n282 1.5005
R485 vdd.n279 vdd.n270 1.5005
R486 vdd.n277 vdd.n276 1.5005
R487 vdd.n275 vdd.n274 1.5005
R488 vdd.n272 vdd.n186 1.5005
R489 vdd.n315 vdd.n185 1.5005
R490 vdd.n318 vdd.n317 1.5005
R491 vdd.n320 vdd.n319 1.5005
R492 vdd.n322 vdd.n321 1.5005
R493 vdd.n184 vdd.n157 1.5005
R494 vdd.n183 vdd.n182 1.5005
R495 vdd.n177 vdd.n176 1.5005
R496 vdd.n175 vdd.n174 1.5005
R497 vdd.n172 vdd.n161 1.5005
R498 vdd.n170 vdd.n169 1.5005
R499 vdd.n168 vdd.n167 1.5005
R500 vdd.n165 vdd.n163 1.5005
R501 vdd.n128 vdd.n127 1.5005
R502 vdd.n335 vdd.n334 1.5005
R503 vdd.n337 vdd.n336 1.5005
R504 vdd.n126 vdd.n109 1.5005
R505 vdd.n125 vdd.n124 1.5005
R506 vdd.n122 vdd.n121 1.5005
R507 vdd.n119 vdd.n111 1.5005
R508 vdd.n117 vdd.n116 1.5005
R509 vdd.n115 vdd.n114 1.5005
R510 vdd.n777 vdd.n9 1.5005
R511 vdd.n776 vdd.n775 1.5005
R512 vdd.n774 vdd.n11 1.5005
R513 vdd.n773 vdd.n772 1.5005
R514 vdd.n771 vdd.n770 1.5005
R515 vdd.n769 vdd.n13 1.5005
R516 vdd.n768 vdd.n767 1.5005
R517 vdd.n762 vdd.n14 1.5005
R518 vdd.n761 vdd.n760 1.5005
R519 vdd.n16 vdd.n15 1.5005
R520 vdd.n740 vdd.n735 1.5005
R521 vdd.n742 vdd.n741 1.5005
R522 vdd.n744 vdd.n734 1.5005
R523 vdd.n746 vdd.n745 1.5005
R524 vdd.n747 vdd.n21 1.5005
R525 vdd.n749 vdd.n748 1.5005
R526 vdd.n733 vdd.n20 1.5005
R527 vdd.n732 vdd.n731 1.5005
R528 vdd.n730 vdd.n22 1.5005
R529 vdd.n729 vdd.n728 1.5005
R530 vdd.n723 vdd.n23 1.5005
R531 vdd.n722 vdd.n721 1.5005
R532 vdd.n719 vdd.n24 1.5005
R533 vdd.n718 vdd.n717 1.5005
R534 vdd.n716 vdd.n25 1.5005
R535 vdd.n714 vdd.n713 1.5005
R536 vdd.n30 vdd.n29 1.5005
R537 vdd.n691 vdd.n690 1.5005
R538 vdd.n693 vdd.n692 1.5005
R539 vdd.n695 vdd.n689 1.5005
R540 vdd.n697 vdd.n696 1.5005
R541 vdd.n699 vdd.n35 1.5005
R542 vdd.n701 vdd.n700 1.5005
R543 vdd.n685 vdd.n34 1.5005
R544 vdd.n684 vdd.n683 1.5005
R545 vdd.n682 vdd.n36 1.5005
R546 vdd.n681 vdd.n680 1.5005
R547 vdd.n678 vdd.n677 1.5005
R548 vdd.n676 vdd.n41 1.5005
R549 vdd.n675 vdd.n674 1.5005
R550 vdd.n673 vdd.n42 1.5005
R551 vdd.n672 vdd.n671 1.5005
R552 vdd.n44 vdd.n43 1.5005
R553 vdd.n647 vdd.n642 1.5005
R554 vdd.n649 vdd.n648 1.5005
R555 vdd.n651 vdd.n641 1.5005
R556 vdd.n653 vdd.n652 1.5005
R557 vdd.n654 vdd.n57 1.5005
R558 vdd.n656 vdd.n655 1.5005
R559 vdd.n639 vdd.n56 1.5005
R560 vdd.n638 vdd.n637 1.5005
R561 vdd.n636 vdd.n61 1.5005
R562 vdd.n635 vdd.n634 1.5005
R563 vdd.n633 vdd.n632 1.5005
R564 vdd.n631 vdd.n63 1.5005
R565 vdd.n630 vdd.n629 1.5005
R566 vdd.n627 vdd.n64 1.5005
R567 vdd.n626 vdd.n625 1.5005
R568 vdd.n69 vdd.n68 1.5005
R569 vdd.n595 vdd.n594 1.5005
R570 vdd.n597 vdd.n596 1.5005
R571 vdd.n598 vdd.n590 1.5005
R572 vdd.n601 vdd.n600 1.5005
R573 vdd.n602 vdd.n589 1.5005
R574 vdd.n604 vdd.n603 1.5005
R575 vdd.n606 vdd.n605 1.5005
R576 vdd.n607 vdd.n587 1.5005
R577 vdd.n609 vdd.n608 1.5005
R578 vdd.n611 vdd.n75 1.5005
R579 vdd.n613 vdd.n612 1.5005
R580 vdd.n583 vdd.n74 1.5005
R581 vdd.n582 vdd.n581 1.5005
R582 vdd.n580 vdd.n76 1.5005
R583 vdd.n579 vdd.n578 1.5005
R584 vdd.n576 vdd.n575 1.5005
R585 vdd.n574 vdd.n81 1.5005
R586 vdd.n573 vdd.n572 1.5005
R587 vdd.n571 vdd.n82 1.5005
R588 vdd.n570 vdd.n569 1.5005
R589 vdd.n84 vdd.n83 1.5005
R590 vdd.n504 vdd.n499 1.5005
R591 vdd.n506 vdd.n505 1.5005
R592 vdd.n508 vdd.n498 1.5005
R593 vdd.n510 vdd.n509 1.5005
R594 vdd.n511 vdd.n493 1.5005
R595 vdd.n513 vdd.n512 1.5005
R596 vdd.n515 vdd.n492 1.5005
R597 vdd.n517 vdd.n516 1.5005
R598 vdd.n518 vdd.n491 1.5005
R599 vdd.n520 vdd.n519 1.5005
R600 vdd.n523 vdd.n490 1.5005
R601 vdd.n525 vdd.n524 1.5005
R602 vdd.n526 vdd.n486 1.5005
R603 vdd.n529 vdd.n528 1.5005
R604 vdd.n531 vdd.n485 1.5005
R605 vdd.n533 vdd.n532 1.5005
R606 vdd.n534 vdd.n368 1.5005
R607 vdd.n536 vdd.n535 1.5005
R608 vdd.n484 vdd.n367 1.5005
R609 vdd.n482 vdd.n481 1.5005
R610 vdd.n480 vdd.n372 1.5005
R611 vdd.n479 vdd.n478 1.5005
R612 vdd.n477 vdd.n476 1.5005
R613 vdd.n475 vdd.n374 1.5005
R614 vdd.n474 vdd.n473 1.5005
R615 vdd.n471 vdd.n375 1.5005
R616 vdd.n470 vdd.n469 1.5005
R617 vdd.n467 vdd.n379 1.5005
R618 vdd.n466 vdd.n465 1.5005
R619 vdd.n464 vdd.n380 1.5005
R620 vdd.n463 vdd.n462 1.5005
R621 vdd.n460 vdd.n459 1.5005
R622 vdd.n458 vdd.n385 1.5005
R623 vdd.n457 vdd.n456 1.5005
R624 vdd.n454 vdd.n386 1.5005
R625 vdd.n453 vdd.n452 1.5005
R626 vdd.n451 vdd.n387 1.5005
R627 vdd.n449 vdd.n448 1.5005
R628 vdd.n446 vdd.n391 1.5005
R629 vdd.n445 vdd.n444 1.5005
R630 vdd.n443 vdd.n392 1.5005
R631 vdd.n442 vdd.n441 1.5005
R632 vdd.n440 vdd.n393 1.5005
R633 vdd.n438 vdd.n437 1.5005
R634 vdd.n432 vdd.n394 1.5005
R635 vdd.n431 vdd.n430 1.5005
R636 vdd.n429 vdd.n395 1.5005
R637 vdd.n427 vdd.n426 1.5005
R638 vdd.n425 vdd.n396 1.5005
R639 vdd.n424 vdd.n423 1.5005
R640 vdd.n422 vdd.n421 1.5005
R641 vdd.n420 vdd.n419 1.5005
R642 vdd.n418 vdd.n402 1.5005
R643 vdd.n417 vdd.n416 1.5005
R644 vdd.n415 vdd.n403 1.5005
R645 vdd.n414 vdd.n413 1.5005
R646 vdd.n268 vdd.n267 1.41716
R647 vdd.n268 vdd.n212 1.37269
R648 vdd.n267 vdd.n213 1.35023
R649 vdd.n263 vdd.n212 1.34472
R650 vdd.n214 vdd.n213 1.2534
R651 vdd.n215 vdd.n214 1.19837
R652 vdd.n324 vdd.n150 1.1005
R653 vdd.n326 vdd.n150 1.1005
R654 vdd.n327 vdd.n141 1.1005
R655 vdd.n327 vdd.n140 1.1005
R656 vdd.n327 vdd.n142 1.1005
R657 vdd.n327 vdd.n139 1.1005
R658 vdd.n327 vdd.n143 1.1005
R659 vdd.n327 vdd.n326 1.1005
R660 vdd.n156 vdd.n136 1.1005
R661 vdd.n156 vdd.n141 1.1005
R662 vdd.n156 vdd.n140 1.1005
R663 vdd.n156 vdd.n142 1.1005
R664 vdd.n156 vdd.n139 1.1005
R665 vdd.n156 vdd.n143 1.1005
R666 vdd.n180 vdd.n156 1.1005
R667 vdd.n324 vdd.n156 1.1005
R668 vdd.n151 vdd.n136 1.1005
R669 vdd.n151 vdd.n141 1.1005
R670 vdd.n151 vdd.n140 1.1005
R671 vdd.n151 vdd.n142 1.1005
R672 vdd.n151 vdd.n139 1.1005
R673 vdd.n151 vdd.n143 1.1005
R674 vdd.n324 vdd.n151 1.1005
R675 vdd.n326 vdd.n151 1.1005
R676 vdd.n154 vdd.n136 1.1005
R677 vdd.n154 vdd.n141 1.1005
R678 vdd.n154 vdd.n140 1.1005
R679 vdd.n154 vdd.n142 1.1005
R680 vdd.n154 vdd.n139 1.1005
R681 vdd.n154 vdd.n143 1.1005
R682 vdd.n324 vdd.n154 1.1005
R683 vdd.n325 vdd.n136 1.1005
R684 vdd.n325 vdd.n141 1.1005
R685 vdd.n325 vdd.n140 1.1005
R686 vdd.n325 vdd.n142 1.1005
R687 vdd.n325 vdd.n139 1.1005
R688 vdd.n325 vdd.n143 1.1005
R689 vdd.n325 vdd.n324 1.1005
R690 vdd.n325 vdd.n153 1.1005
R691 vdd.n326 vdd.n325 1.1005
R692 vdd.n345 vdd.n105 1.1005
R693 vdd.n345 vdd.n93 1.1005
R694 vdd.n345 vdd.n92 1.1005
R695 vdd.n343 vdd.n92 1.1005
R696 vdd.n105 vdd.n103 1.1005
R697 vdd.n103 vdd.n95 1.1005
R698 vdd.n103 vdd.n97 1.1005
R699 vdd.n103 vdd.n94 1.1005
R700 vdd.n350 vdd.n103 1.1005
R701 vdd.n103 vdd.n93 1.1005
R702 vdd.n103 vdd.n92 1.1005
R703 vdd.n105 vdd.n100 1.1005
R704 vdd.n100 vdd.n95 1.1005
R705 vdd.n100 vdd.n97 1.1005
R706 vdd.n100 vdd.n94 1.1005
R707 vdd.n350 vdd.n100 1.1005
R708 vdd.n100 vdd.n93 1.1005
R709 vdd.n100 vdd.n92 1.1005
R710 vdd.n349 vdd.n105 1.1005
R711 vdd.n349 vdd.n95 1.1005
R712 vdd.n349 vdd.n97 1.1005
R713 vdd.n349 vdd.n94 1.1005
R714 vdd.n350 vdd.n349 1.1005
R715 vdd.n349 vdd.n93 1.1005
R716 vdd.n349 vdd.n92 1.1005
R717 vdd.n105 vdd.n99 1.1005
R718 vdd.n99 vdd.n95 1.1005
R719 vdd.n99 vdd.n97 1.1005
R720 vdd.n99 vdd.n94 1.1005
R721 vdd.n350 vdd.n99 1.1005
R722 vdd.n99 vdd.n92 1.1005
R723 vdd.n351 vdd.n95 1.1005
R724 vdd.n351 vdd.n97 1.1005
R725 vdd.n351 vdd.n94 1.1005
R726 vdd.n351 vdd.n350 1.1005
R727 vdd.n351 vdd.n93 1.1005
R728 vdd.n351 vdd.n92 1.1005
R729 vdd.n557 vdd.n88 1.1005
R730 vdd.n559 vdd.n558 1.1005
R731 vdd.n560 vdd.n48 1.1005
R732 vdd.n662 vdd.n661 1.1005
R733 vdd.n663 vdd.n47 1.1005
R734 vdd.n665 vdd.n664 1.1005
R735 vdd.n667 vdd.n1 1.1005
R736 vdd.n784 vdd.n2 1.1005
R737 vdd.n207 vdd.n193 1.1005
R738 vdd.n207 vdd.n194 1.1005
R739 vdd.n310 vdd.n207 1.1005
R740 vdd.n201 vdd.n187 1.1005
R741 vdd.n201 vdd.n194 1.1005
R742 vdd.n310 vdd.n201 1.1005
R743 vdd.n311 vdd.n187 1.1005
R744 vdd.n311 vdd.n191 1.1005
R745 vdd.n311 vdd.n192 1.1005
R746 vdd.n311 vdd.n190 1.1005
R747 vdd.n311 vdd.n193 1.1005
R748 vdd.n311 vdd.n194 1.1005
R749 vdd.n311 vdd.n310 1.1005
R750 vdd.n198 vdd.n187 1.1005
R751 vdd.n198 vdd.n191 1.1005
R752 vdd.n198 vdd.n192 1.1005
R753 vdd.n198 vdd.n190 1.1005
R754 vdd.n198 vdd.n193 1.1005
R755 vdd.n198 vdd.n194 1.1005
R756 vdd.n310 vdd.n198 1.1005
R757 vdd.n309 vdd.n187 1.1005
R758 vdd.n309 vdd.n191 1.1005
R759 vdd.n309 vdd.n192 1.1005
R760 vdd.n309 vdd.n190 1.1005
R761 vdd.n309 vdd.n193 1.1005
R762 vdd.n309 vdd.n194 1.1005
R763 vdd.n310 vdd.n309 1.1005
R764 vdd.n197 vdd.n187 1.1005
R765 vdd.n197 vdd.n191 1.1005
R766 vdd.n197 vdd.n192 1.1005
R767 vdd.n197 vdd.n190 1.1005
R768 vdd.n197 vdd.n194 1.1005
R769 vdd.n310 vdd.n197 1.1005
R770 vdd.n187 vdd.n0 1.1005
R771 vdd.n191 vdd.n0 1.1005
R772 vdd.n192 vdd.n0 1.1005
R773 vdd.n190 vdd.n0 1.1005
R774 vdd.n193 vdd.n0 1.1005
R775 vdd.n310 vdd.n0 1.1005
R776 vdd.n783 vdd.n782 1.1005
R777 vdd.n407 vdd 0.83073
R778 vdd.n400 vdd 0.83073
R779 vdd.n436 vdd 0.83073
R780 vdd.n450 vdd 0.83073
R781 vdd.n384 vdd 0.83073
R782 vdd.n472 vdd 0.83073
R783 vdd.n483 vdd 0.83073
R784 vdd.n527 vdd 0.83073
R785 vdd.n497 vdd 0.83073
R786 vdd.n503 vdd 0.83073
R787 vdd.n577 vdd 0.83073
R788 vdd.n610 vdd 0.83073
R789 vdd.n599 vdd 0.83073
R790 vdd.n628 vdd 0.83073
R791 vdd.n640 vdd 0.83073
R792 vdd.n646 vdd 0.83073
R793 vdd.n679 vdd 0.83073
R794 vdd.n698 vdd 0.83073
R795 vdd.n715 vdd 0.83073
R796 vdd.n727 vdd 0.83073
R797 vdd.n739 vdd 0.83073
R798 vdd.n766 vdd 0.83073
R799 vdd.n269 vdd.n268 0.765466
R800 vdd.n779 vdd.n778 0.762052
R801 vdd.n405 vdd.n404 0.698729
R802 vdd.n406 vdd.n405 0.698729
R803 vdd.n398 vdd.n397 0.698729
R804 vdd.n399 vdd.n398 0.698729
R805 vdd.n434 vdd.n433 0.698729
R806 vdd.n435 vdd.n434 0.698729
R807 vdd.n389 vdd.n388 0.698729
R808 vdd.n390 vdd.n389 0.698729
R809 vdd.n382 vdd.n381 0.698729
R810 vdd.n383 vdd.n382 0.698729
R811 vdd.n377 vdd.n376 0.698729
R812 vdd.n378 vdd.n377 0.698729
R813 vdd.n370 vdd.n369 0.698729
R814 vdd.n371 vdd.n370 0.698729
R815 vdd.n488 vdd.n487 0.698729
R816 vdd.n489 vdd.n488 0.698729
R817 vdd.n495 vdd.n494 0.698729
R818 vdd.n496 vdd.n495 0.698729
R819 vdd.n501 vdd.n500 0.698729
R820 vdd.n502 vdd.n501 0.698729
R821 vdd.n79 vdd.n78 0.698729
R822 vdd.n80 vdd.n79 0.698729
R823 vdd.n585 vdd.n584 0.698729
R824 vdd.n586 vdd.n585 0.698729
R825 vdd.n592 vdd.n591 0.698729
R826 vdd.n593 vdd.n592 0.698729
R827 vdd.n66 vdd.n65 0.698729
R828 vdd.n67 vdd.n66 0.698729
R829 vdd.n59 vdd.n58 0.698729
R830 vdd.n60 vdd.n59 0.698729
R831 vdd.n644 vdd.n643 0.698729
R832 vdd.n645 vdd.n644 0.698729
R833 vdd.n39 vdd.n38 0.698729
R834 vdd.n40 vdd.n39 0.698729
R835 vdd.n687 vdd.n686 0.698729
R836 vdd.n688 vdd.n687 0.698729
R837 vdd.n27 vdd.n26 0.698729
R838 vdd.n28 vdd.n27 0.698729
R839 vdd.n725 vdd.n724 0.698729
R840 vdd.n726 vdd.n725 0.698729
R841 vdd.n737 vdd.n736 0.698729
R842 vdd.n738 vdd.n737 0.698729
R843 vdd.n764 vdd.n763 0.698729
R844 vdd.n765 vdd.n764 0.698729
R845 vdd.n288 vdd 0.6957
R846 vdd.n153 vdd.n137 0.5507
R847 vdd.n328 vdd.n136 0.5507
R848 vdd.n326 vdd.n131 0.5507
R849 vdd.n155 vdd.n153 0.5507
R850 vdd.n180 vdd.n179 0.5507
R851 vdd.n180 vdd.n152 0.5507
R852 vdd.n347 vdd.n346 0.5507
R853 vdd.n340 vdd.n339 0.5507
R854 vdd.n347 vdd.n107 0.5507
R855 vdd.n339 vdd.n104 0.5507
R856 vdd.n348 vdd.n347 0.5507
R857 vdd.n339 vdd.n91 0.5507
R858 vdd.n204 vdd.n196 0.5507
R859 vdd.n307 vdd.n189 0.5507
R860 vdd.n196 vdd.n188 0.5507
R861 vdd.n308 vdd.n307 0.5507
R862 vdd.n208 vdd.n196 0.5507
R863 vdd.n307 vdd.n306 0.5507
R864 vdd.n150 vdd.n149 0.5505
R865 vdd.n150 vdd.n148 0.5505
R866 vdd.n150 vdd.n147 0.5505
R867 vdd.n327 vdd.n138 0.5505
R868 vdd.n329 vdd.n135 0.5505
R869 vdd.n329 vdd.n134 0.5505
R870 vdd.n329 vdd.n133 0.5505
R871 vdd.n329 vdd.n132 0.5505
R872 vdd.n154 vdd.n144 0.5505
R873 vdd.n345 vdd.n344 0.5505
R874 vdd.n345 vdd.n98 0.5505
R875 vdd.n343 vdd.n342 0.5505
R876 vdd.n343 vdd.n341 0.5505
R877 vdd.n343 vdd.n102 0.5505
R878 vdd.n108 vdd.n99 0.5505
R879 vdd.n351 vdd.n96 0.5505
R880 vdd.n207 vdd.n206 0.5505
R881 vdd.n207 vdd.n205 0.5505
R882 vdd.n201 vdd.n200 0.5505
R883 vdd.n201 vdd.n199 0.5505
R884 vdd.n209 vdd.n197 0.5505
R885 vdd.n195 vdd.n0 0.5505
R886 vdd.n556 vdd.n90 0.549388
R887 vdd.n556 vdd.n555 0.548016
R888 vdd.n556 vdd.n354 0.548016
R889 vdd.n556 vdd.n353 0.548016
R890 vdd.n556 vdd.n352 0.548016
R891 vdd.n662 vdd.n49 0.548016
R892 vdd.n662 vdd.n50 0.548016
R893 vdd.n662 vdd.n51 0.548016
R894 vdd.n662 vdd.n52 0.548016
R895 vdd.n784 vdd.n6 0.548016
R896 vdd.n784 vdd.n5 0.548016
R897 vdd.n784 vdd.n4 0.548016
R898 vdd.n784 vdd.n3 0.548016
R899 vdd.n223 vdd.n222 0.328961
R900 vdd.n257 vdd.n256 0.328961
R901 vdd.n115 vdd.n106 0.325781
R902 vdd.n408 vdd.n407 0.323766
R903 vdd.n236 vdd.n235 0.322808
R904 vdd.n245 vdd.n244 0.322188
R905 vdd vdd.n406 0.317156
R906 vdd vdd.n399 0.317156
R907 vdd vdd.n435 0.317156
R908 vdd vdd.n390 0.317156
R909 vdd vdd.n383 0.317156
R910 vdd vdd.n378 0.317156
R911 vdd vdd.n371 0.317156
R912 vdd vdd.n489 0.317156
R913 vdd vdd.n496 0.317156
R914 vdd vdd.n502 0.317156
R915 vdd vdd.n80 0.317156
R916 vdd vdd.n586 0.317156
R917 vdd vdd.n593 0.317156
R918 vdd vdd.n67 0.317156
R919 vdd vdd.n60 0.317156
R920 vdd vdd.n645 0.317156
R921 vdd vdd.n40 0.317156
R922 vdd vdd.n688 0.317156
R923 vdd vdd.n28 0.317156
R924 vdd vdd.n726 0.317156
R925 vdd vdd.n738 0.317156
R926 vdd vdd.n765 0.317156
R927 vdd.n292 vdd.n291 0.316786
R928 vdd.n248 vdd.n247 0.316029
R929 vdd.n233 vdd.n232 0.31602
R930 vdd.n293 vdd.n292 0.314786
R931 vdd.n295 vdd.n203 0.314786
R932 vdd.n310 vdd.n202 0.314786
R933 vdd.n300 vdd.n196 0.314786
R934 vdd.n211 vdd.n194 0.314786
R935 vdd.n307 vdd.n305 0.314786
R936 vdd.n281 vdd.n193 0.314786
R937 vdd.n280 vdd.n190 0.314786
R938 vdd.n278 vdd.n192 0.314786
R939 vdd.n271 vdd.n191 0.314786
R940 vdd.n273 vdd.n187 0.314786
R941 vdd.n314 vdd.n313 0.314786
R942 vdd.n316 vdd.n146 0.314786
R943 vdd.n326 vdd.n145 0.314786
R944 vdd.n158 vdd.n153 0.314786
R945 vdd.n324 vdd.n323 0.314786
R946 vdd.n181 vdd.n180 0.314786
R947 vdd.n178 vdd.n143 0.314786
R948 vdd.n160 vdd.n139 0.314786
R949 vdd.n173 vdd.n142 0.314786
R950 vdd.n171 vdd.n140 0.314786
R951 vdd.n162 vdd.n141 0.314786
R952 vdd.n166 vdd.n136 0.314786
R953 vdd.n164 vdd.n129 0.314786
R954 vdd.n333 vdd.n332 0.314786
R955 vdd.n110 vdd.n92 0.314786
R956 vdd.n339 vdd.n338 0.314786
R957 vdd.n123 vdd.n93 0.314786
R958 vdd.n350 vdd.n101 0.314786
R959 vdd.n120 vdd.n94 0.314786
R960 vdd.n118 vdd.n97 0.314786
R961 vdd.n112 vdd.n95 0.314786
R962 vdd.n113 vdd.n105 0.314786
R963 vdd.n260 vdd.n259 0.309867
R964 vdd.n226 vdd.n225 0.309867
R965 vdd.n255 vdd.n254 0.309247
R966 vdd.n221 vdd.n220 0.309247
R967 vdd.n238 vdd.n237 0.303088
R968 vdd.n243 vdd.n242 0.303079
R969 vdd.n250 vdd.n249 0.296926
R970 vdd.n216 vdd.n215 0.296926
R971 vdd.n265 vdd.n263 0.296305
R972 vdd.n231 vdd.n230 0.296305
R973 vdd.n225 vdd.n224 0.291089
R974 vdd.n259 vdd.n258 0.291089
R975 vdd.n262 vdd.n261 0.290146
R976 vdd.n228 vdd.n227 0.290146
R977 vdd.n219 vdd.n218 0.290137
R978 vdd.n253 vdd.n252 0.290137
R979 vdd.n234 vdd.n233 0.284975
R980 vdd.n247 vdd.n246 0.284443
R981 vdd.n240 vdd.n239 0.283985
R982 vdd.n241 vdd.n240 0.283364
R983 vdd.n246 vdd.n245 0.278673
R984 vdd.n235 vdd.n234 0.278148
R985 vdd.n252 vdd.n251 0.277205
R986 vdd.n218 vdd.n217 0.277205
R987 vdd.n229 vdd.n228 0.277196
R988 vdd.n264 vdd.n262 0.277196
R989 vdd.n224 vdd.n223 0.272034
R990 vdd.n258 vdd.n257 0.272034
R991 vdd.n265 vdd.n264 0.271044
R992 vdd.n230 vdd.n229 0.271044
R993 vdd.n251 vdd.n250 0.270423
R994 vdd.n217 vdd.n216 0.270423
R995 vdd.n242 vdd.n241 0.264264
R996 vdd.n239 vdd.n238 0.264255
R997 vdd.n254 vdd.n253 0.258102
R998 vdd.n220 vdd.n219 0.258102
R999 vdd.n261 vdd.n260 0.257482
R1000 vdd.n227 vdd.n226 0.257482
R1001 vdd.n232 vdd.n231 0.251323
R1002 vdd.n249 vdd.n248 0.251314
R1003 vdd.n556 vdd 0.248
R1004 vdd.n244 vdd.n243 0.245161
R1005 vdd.n237 vdd.n236 0.244541
R1006 vdd.n256 vdd.n255 0.238382
R1007 vdd.n222 vdd.n221 0.238382
R1008 vdd.n159 vdd 0.217715
R1009 vdd.n266 vdd.n214 0.166751
R1010 vdd.n662 vdd 0.16242
R1011 vdd.n332 vdd.n331 0.157643
R1012 vdd.n330 vdd.n129 0.157643
R1013 vdd.n146 vdd.n130 0.157643
R1014 vdd.n313 vdd.n312 0.157643
R1015 vdd.n10 vdd 0.119054
R1016 vdd.n270 vdd.n269 0.100015
R1017 vdd.n269 vdd 0.096503
R1018 vdd.n662 vdd 0.0845153
R1019 vdd.n556 vdd 0.0845153
R1020 vdd vdd.n784 0.0845153
R1021 vdd.n347 vdd.n106 0.0840543
R1022 vdd.n784 vdd 0.0768767
R1023 vdd.n411 vdd.n410 0.0591667
R1024 vdd.n411 vdd.n358 0.0591667
R1025 vdd.n359 vdd.n358 0.0591667
R1026 vdd.n360 vdd.n359 0.0591667
R1027 vdd.n361 vdd.n360 0.0591667
R1028 vdd.n362 vdd.n361 0.0591667
R1029 vdd.n363 vdd.n362 0.0591667
R1030 vdd.n364 vdd.n363 0.0591667
R1031 vdd.n365 vdd.n364 0.0591667
R1032 vdd.n538 vdd.n365 0.0591667
R1033 vdd.n538 vdd.n366 0.0591667
R1034 vdd.n521 vdd.n366 0.0591667
R1035 vdd.n521 vdd.n87 0.0591667
R1036 vdd.n87 vdd.n85 0.0591667
R1037 vdd.n567 vdd.n85 0.0591667
R1038 vdd.n567 vdd.n73 0.0591667
R1039 vdd.n614 vdd.n73 0.0591667
R1040 vdd.n614 vdd.n70 0.0591667
R1041 vdd.n622 vdd.n70 0.0591667
R1042 vdd.n623 vdd.n622 0.0591667
R1043 vdd.n623 vdd.n55 0.0591667
R1044 vdd.n658 vdd.n55 0.0591667
R1045 vdd.n658 vdd.n45 0.0591667
R1046 vdd.n669 vdd.n45 0.0591667
R1047 vdd.n669 vdd.n33 0.0591667
R1048 vdd.n703 vdd.n33 0.0591667
R1049 vdd.n703 vdd.n31 0.0591667
R1050 vdd.n711 vdd.n31 0.0591667
R1051 vdd.n711 vdd.n19 0.0591667
R1052 vdd.n751 vdd.n19 0.0591667
R1053 vdd.n751 vdd.n17 0.0591667
R1054 vdd.n758 vdd.n17 0.0591667
R1055 vdd.n758 vdd.n8 0.0591667
R1056 vdd.n780 vdd.n8 0.0591667
R1057 vdd.n409 vdd.n357 0.0591667
R1058 vdd.n553 vdd.n357 0.0591667
R1059 vdd.n553 vdd.n552 0.0591667
R1060 vdd.n552 vdd.n551 0.0591667
R1061 vdd.n551 vdd.n549 0.0591667
R1062 vdd.n549 vdd.n546 0.0591667
R1063 vdd.n546 vdd.n545 0.0591667
R1064 vdd.n545 vdd.n542 0.0591667
R1065 vdd.n542 vdd.n541 0.0591667
R1066 vdd.n541 vdd.n539 0.0591667
R1067 vdd.n539 vdd.n89 0.0591667
R1068 vdd.n89 vdd.n86 0.0591667
R1069 vdd.n562 vdd.n86 0.0591667
R1070 vdd.n563 vdd.n562 0.0591667
R1071 vdd.n566 vdd.n563 0.0591667
R1072 vdd.n566 vdd.n72 0.0591667
R1073 vdd.n617 vdd.n72 0.0591667
R1074 vdd.n618 vdd.n617 0.0591667
R1075 vdd.n621 vdd.n618 0.0591667
R1076 vdd.n621 vdd.n54 0.0591667
R1077 vdd.n660 vdd.n54 0.0591667
R1078 vdd.n660 vdd.n659 0.0591667
R1079 vdd.n659 vdd.n46 0.0591667
R1080 vdd.n668 vdd.n46 0.0591667
R1081 vdd.n668 vdd.n32 0.0591667
R1082 vdd.n704 vdd.n32 0.0591667
R1083 vdd.n707 vdd.n704 0.0591667
R1084 vdd.n710 vdd.n707 0.0591667
R1085 vdd.n710 vdd.n18 0.0591667
R1086 vdd.n752 vdd.n18 0.0591667
R1087 vdd.n755 vdd.n752 0.0591667
R1088 vdd.n757 vdd.n755 0.0591667
R1089 vdd.n757 vdd.n7 0.0591667
R1090 vdd.n781 vdd.n7 0.0591667
R1091 vdd.n213 vdd 0.0555
R1092 vdd.n266 vdd.t0 0.0507959
R1093 vdd.n413 vdd.n408 0.0374917
R1094 vdd.n329 vdd 0.0310507
R1095 vdd.n778 vdd.n777 0.02024
R1096 vdd.n113 vdd.n106 0.0183783
R1097 vdd.n415 vdd.n414 0.0148733
R1098 vdd.n416 vdd.n415 0.0148733
R1099 vdd.n416 vdd.n402 0.0148733
R1100 vdd.n420 vdd.n402 0.0148733
R1101 vdd.n421 vdd.n420 0.0148733
R1102 vdd.n425 vdd.n424 0.0148733
R1103 vdd.n426 vdd.n425 0.0148733
R1104 vdd.n426 vdd.n395 0.0148733
R1105 vdd.n431 vdd.n395 0.0148733
R1106 vdd.n432 vdd.n431 0.0148733
R1107 vdd.n437 vdd.n432 0.0148733
R1108 vdd.n442 vdd.n393 0.0148733
R1109 vdd.n443 vdd.n442 0.0148733
R1110 vdd.n444 vdd.n443 0.0148733
R1111 vdd.n444 vdd.n391 0.0148733
R1112 vdd.n449 vdd.n391 0.0148733
R1113 vdd.n452 vdd.n451 0.0148733
R1114 vdd.n452 vdd.n386 0.0148733
R1115 vdd.n457 vdd.n386 0.0148733
R1116 vdd.n458 vdd.n457 0.0148733
R1117 vdd.n459 vdd.n458 0.0148733
R1118 vdd.n464 vdd.n463 0.0148733
R1119 vdd.n465 vdd.n464 0.0148733
R1120 vdd.n465 vdd.n379 0.0148733
R1121 vdd.n470 vdd.n379 0.0148733
R1122 vdd.n471 vdd.n470 0.0148733
R1123 vdd.n473 vdd.n374 0.0148733
R1124 vdd.n477 vdd.n374 0.0148733
R1125 vdd.n478 vdd.n477 0.0148733
R1126 vdd.n478 vdd.n372 0.0148733
R1127 vdd.n482 vdd.n372 0.0148733
R1128 vdd.n535 vdd.n484 0.0148733
R1129 vdd.n535 vdd.n534 0.0148733
R1130 vdd.n534 vdd.n533 0.0148733
R1131 vdd.n533 vdd.n485 0.0148733
R1132 vdd.n528 vdd.n485 0.0148733
R1133 vdd.n526 vdd.n525 0.0148733
R1134 vdd.n525 vdd.n490 0.0148733
R1135 vdd.n519 vdd.n490 0.0148733
R1136 vdd.n519 vdd.n518 0.0148733
R1137 vdd.n518 vdd.n517 0.0148733
R1138 vdd.n517 vdd.n492 0.0148733
R1139 vdd.n512 vdd.n511 0.0148733
R1140 vdd.n511 vdd.n510 0.0148733
R1141 vdd.n510 vdd.n498 0.0148733
R1142 vdd.n505 vdd.n498 0.0148733
R1143 vdd.n505 vdd.n504 0.0148733
R1144 vdd.n570 vdd.n83 0.0148733
R1145 vdd.n571 vdd.n570 0.0148733
R1146 vdd.n572 vdd.n571 0.0148733
R1147 vdd.n572 vdd.n81 0.0148733
R1148 vdd.n576 vdd.n81 0.0148733
R1149 vdd.n578 vdd.n76 0.0148733
R1150 vdd.n582 vdd.n76 0.0148733
R1151 vdd.n583 vdd.n582 0.0148733
R1152 vdd.n612 vdd.n583 0.0148733
R1153 vdd.n612 vdd.n611 0.0148733
R1154 vdd.n609 vdd.n587 0.0148733
R1155 vdd.n605 vdd.n587 0.0148733
R1156 vdd.n605 vdd.n604 0.0148733
R1157 vdd.n604 vdd.n589 0.0148733
R1158 vdd.n600 vdd.n589 0.0148733
R1159 vdd.n598 vdd.n597 0.0148733
R1160 vdd.n597 vdd.n594 0.0148733
R1161 vdd.n594 vdd.n68 0.0148733
R1162 vdd.n626 vdd.n68 0.0148733
R1163 vdd.n627 vdd.n626 0.0148733
R1164 vdd.n629 vdd.n63 0.0148733
R1165 vdd.n633 vdd.n63 0.0148733
R1166 vdd.n634 vdd.n633 0.0148733
R1167 vdd.n634 vdd.n61 0.0148733
R1168 vdd.n638 vdd.n61 0.0148733
R1169 vdd.n639 vdd.n638 0.0148733
R1170 vdd.n655 vdd.n654 0.0148733
R1171 vdd.n654 vdd.n653 0.0148733
R1172 vdd.n653 vdd.n641 0.0148733
R1173 vdd.n648 vdd.n641 0.0148733
R1174 vdd.n648 vdd.n647 0.0148733
R1175 vdd.n672 vdd.n43 0.0148733
R1176 vdd.n673 vdd.n672 0.0148733
R1177 vdd.n674 vdd.n673 0.0148733
R1178 vdd.n674 vdd.n41 0.0148733
R1179 vdd.n678 vdd.n41 0.0148733
R1180 vdd.n680 vdd.n36 0.0148733
R1181 vdd.n684 vdd.n36 0.0148733
R1182 vdd.n685 vdd.n684 0.0148733
R1183 vdd.n700 vdd.n685 0.0148733
R1184 vdd.n700 vdd.n699 0.0148733
R1185 vdd.n697 vdd.n689 0.0148733
R1186 vdd.n692 vdd.n689 0.0148733
R1187 vdd.n692 vdd.n691 0.0148733
R1188 vdd.n691 vdd.n29 0.0148733
R1189 vdd.n714 vdd.n29 0.0148733
R1190 vdd.n717 vdd.n716 0.0148733
R1191 vdd.n717 vdd.n24 0.0148733
R1192 vdd.n722 vdd.n24 0.0148733
R1193 vdd.n723 vdd.n722 0.0148733
R1194 vdd.n728 vdd.n723 0.0148733
R1195 vdd.n732 vdd.n22 0.0148733
R1196 vdd.n733 vdd.n732 0.0148733
R1197 vdd.n748 vdd.n733 0.0148733
R1198 vdd.n748 vdd.n747 0.0148733
R1199 vdd.n747 vdd.n746 0.0148733
R1200 vdd.n746 vdd.n734 0.0148733
R1201 vdd.n741 vdd.n740 0.0148733
R1202 vdd.n740 vdd.n15 0.0148733
R1203 vdd.n761 vdd.n15 0.0148733
R1204 vdd.n762 vdd.n761 0.0148733
R1205 vdd.n767 vdd.n762 0.0148733
R1206 vdd.n771 vdd.n13 0.0148733
R1207 vdd.n772 vdd.n771 0.0148733
R1208 vdd.n772 vdd.n11 0.0148733
R1209 vdd.n776 vdd.n11 0.0148733
R1210 vdd.n777 vdd.n776 0.0148733
R1211 vdd.n417 vdd.n403 0.0148733
R1212 vdd.n418 vdd.n417 0.0148733
R1213 vdd.n419 vdd.n418 0.0148733
R1214 vdd.n423 vdd.n422 0.0148733
R1215 vdd.n423 vdd.n396 0.0148733
R1216 vdd.n427 vdd.n396 0.0148733
R1217 vdd.n430 vdd.n429 0.0148733
R1218 vdd.n430 vdd.n394 0.0148733
R1219 vdd.n438 vdd.n394 0.0148733
R1220 vdd.n441 vdd.n440 0.0148733
R1221 vdd.n441 vdd.n392 0.0148733
R1222 vdd.n445 vdd.n392 0.0148733
R1223 vdd.n446 vdd.n445 0.0148733
R1224 vdd.n448 vdd.n387 0.0148733
R1225 vdd.n453 vdd.n387 0.0148733
R1226 vdd.n454 vdd.n453 0.0148733
R1227 vdd.n456 vdd.n385 0.0148733
R1228 vdd.n460 vdd.n385 0.0148733
R1229 vdd.n462 vdd.n460 0.0148733
R1230 vdd.n466 vdd.n380 0.0148733
R1231 vdd.n467 vdd.n466 0.0148733
R1232 vdd.n469 vdd.n467 0.0148733
R1233 vdd.n474 vdd.n375 0.0148733
R1234 vdd.n475 vdd.n474 0.0148733
R1235 vdd.n476 vdd.n475 0.0148733
R1236 vdd.n480 vdd.n479 0.0148733
R1237 vdd.n481 vdd.n480 0.0148733
R1238 vdd.n481 vdd.n367 0.0148733
R1239 vdd.n536 vdd.n368 0.0148733
R1240 vdd.n532 vdd.n368 0.0148733
R1241 vdd.n532 vdd.n531 0.0148733
R1242 vdd.n529 vdd.n486 0.0148733
R1243 vdd.n524 vdd.n486 0.0148733
R1244 vdd.n524 vdd.n523 0.0148733
R1245 vdd.n520 vdd.n491 0.0148733
R1246 vdd.n516 vdd.n491 0.0148733
R1247 vdd.n516 vdd.n515 0.0148733
R1248 vdd.n513 vdd.n493 0.0148733
R1249 vdd.n509 vdd.n493 0.0148733
R1250 vdd.n509 vdd.n508 0.0148733
R1251 vdd.n506 vdd.n499 0.0148733
R1252 vdd.n499 vdd.n84 0.0148733
R1253 vdd.n569 vdd.n84 0.0148733
R1254 vdd.n573 vdd.n82 0.0148733
R1255 vdd.n574 vdd.n573 0.0148733
R1256 vdd.n575 vdd.n574 0.0148733
R1257 vdd.n580 vdd.n579 0.0148733
R1258 vdd.n581 vdd.n580 0.0148733
R1259 vdd.n581 vdd.n74 0.0148733
R1260 vdd.n613 vdd.n74 0.0148733
R1261 vdd.n613 vdd.n75 0.0148733
R1262 vdd.n608 vdd.n75 0.0148733
R1263 vdd.n608 vdd.n607 0.0148733
R1264 vdd.n607 vdd.n606 0.0148733
R1265 vdd.n603 vdd.n602 0.0148733
R1266 vdd.n602 vdd.n601 0.0148733
R1267 vdd.n601 vdd.n590 0.0148733
R1268 vdd.n596 vdd.n595 0.0148733
R1269 vdd.n595 vdd.n69 0.0148733
R1270 vdd.n625 vdd.n69 0.0148733
R1271 vdd.n630 vdd.n64 0.0148733
R1272 vdd.n631 vdd.n630 0.0148733
R1273 vdd.n632 vdd.n631 0.0148733
R1274 vdd.n636 vdd.n635 0.0148733
R1275 vdd.n637 vdd.n636 0.0148733
R1276 vdd.n637 vdd.n56 0.0148733
R1277 vdd.n656 vdd.n57 0.0148733
R1278 vdd.n652 vdd.n57 0.0148733
R1279 vdd.n652 vdd.n651 0.0148733
R1280 vdd.n649 vdd.n642 0.0148733
R1281 vdd.n642 vdd.n44 0.0148733
R1282 vdd.n671 vdd.n44 0.0148733
R1283 vdd.n675 vdd.n42 0.0148733
R1284 vdd.n676 vdd.n675 0.0148733
R1285 vdd.n677 vdd.n676 0.0148733
R1286 vdd.n682 vdd.n681 0.0148733
R1287 vdd.n683 vdd.n682 0.0148733
R1288 vdd.n683 vdd.n34 0.0148733
R1289 vdd.n701 vdd.n35 0.0148733
R1290 vdd.n696 vdd.n35 0.0148733
R1291 vdd.n696 vdd.n695 0.0148733
R1292 vdd.n693 vdd.n690 0.0148733
R1293 vdd.n690 vdd.n30 0.0148733
R1294 vdd.n713 vdd.n30 0.0148733
R1295 vdd.n718 vdd.n25 0.0148733
R1296 vdd.n719 vdd.n718 0.0148733
R1297 vdd.n721 vdd.n719 0.0148733
R1298 vdd.n729 vdd.n23 0.0148733
R1299 vdd.n730 vdd.n729 0.0148733
R1300 vdd.n731 vdd.n730 0.0148733
R1301 vdd.n731 vdd.n20 0.0148733
R1302 vdd.n749 vdd.n21 0.0148733
R1303 vdd.n745 vdd.n21 0.0148733
R1304 vdd.n745 vdd.n744 0.0148733
R1305 vdd.n742 vdd.n735 0.0148733
R1306 vdd.n735 vdd.n16 0.0148733
R1307 vdd.n760 vdd.n16 0.0148733
R1308 vdd.n768 vdd.n14 0.0148733
R1309 vdd.n769 vdd.n768 0.0148733
R1310 vdd.n770 vdd.n769 0.0148733
R1311 vdd.n774 vdd.n773 0.0148733
R1312 vdd.n775 vdd.n774 0.0148733
R1313 vdd.n775 vdd.n9 0.0148733
R1314 vdd.n741 vdd.n739 0.0147267
R1315 vdd.n448 vdd.n447 0.01458
R1316 vdd.n721 vdd.n720 0.01458
R1317 vdd.n655 vdd.n640 0.0144333
R1318 vdd.n267 vdd.n266 0.0142662
R1319 vdd.n512 vdd.n497 0.01414
R1320 vdd.n439 vdd.n438 0.0139933
R1321 vdd.n750 vdd.n749 0.0139933
R1322 vdd.n311 vdd 0.013942
R1323 vdd.n436 vdd.n393 0.0138467
R1324 vdd.n575 vdd.n77 0.0137
R1325 vdd.n603 vdd.n588 0.0137
R1326 vdd.n421 vdd.n400 0.0135533
R1327 vdd.n456 vdd.n455 0.0134067
R1328 vdd.n713 vdd.n712 0.0134067
R1329 vdd.n528 vdd.n527 0.01326
R1330 vdd.n628 vdd.n627 0.0129667
R1331 vdd.n428 vdd.n427 0.01282
R1332 vdd.n743 vdd.n742 0.01282
R1333 vdd.n728 vdd.n727 0.0126733
R1334 vdd.n569 vdd.n568 0.0125267
R1335 vdd.n596 vdd.n71 0.0125267
R1336 vdd.n554 vdd.n356 0.0125
R1337 vdd.n550 vdd.n355 0.0125
R1338 vdd.n548 vdd.n547 0.0125
R1339 vdd.n544 vdd.n543 0.0125
R1340 vdd.n540 vdd.n88 0.0125
R1341 vdd.n559 vdd.n88 0.0125
R1342 vdd.n560 vdd.n559 0.0125
R1343 vdd.n561 vdd.n560 0.0125
R1344 vdd.n565 vdd.n564 0.0125
R1345 vdd.n616 vdd.n615 0.0125
R1346 vdd.n620 vdd.n619 0.0125
R1347 vdd.n661 vdd.n53 0.0125
R1348 vdd.n661 vdd.n47 0.0125
R1349 vdd.n665 vdd.n47 0.0125
R1350 vdd.n667 vdd.n665 0.0125
R1351 vdd.n667 vdd.n666 0.0125
R1352 vdd.n706 vdd.n705 0.0125
R1353 vdd.n709 vdd.n708 0.0125
R1354 vdd.n754 vdd.n753 0.0125
R1355 vdd.n756 vdd.n2 0.0125
R1356 vdd.n782 vdd.n2 0.0125
R1357 vdd.n766 vdd.n13 0.01238
R1358 vdd.n461 vdd.n380 0.0122333
R1359 vdd.n695 vdd.n694 0.0122333
R1360 vdd.n646 vdd.n43 0.0120867
R1361 vdd.n503 vdd.n83 0.0117933
R1362 vdd.n419 vdd.n401 0.0116467
R1363 vdd.n759 vdd.n14 0.0116467
R1364 vdd.n116 vdd.n115 0.0116392
R1365 vdd.n116 vdd.n111 0.0116392
R1366 vdd.n122 vdd.n111 0.0116392
R1367 vdd.n125 vdd.n122 0.0116392
R1368 vdd.n126 vdd.n125 0.0116392
R1369 vdd.n336 vdd.n126 0.0116392
R1370 vdd.n336 vdd.n335 0.0116392
R1371 vdd.n335 vdd.n127 0.0116392
R1372 vdd.n163 vdd.n127 0.0116392
R1373 vdd.n168 vdd.n163 0.0116392
R1374 vdd.n169 vdd.n168 0.0116392
R1375 vdd.n169 vdd.n161 0.0116392
R1376 vdd.n175 vdd.n161 0.0116392
R1377 vdd.n176 vdd.n175 0.0116392
R1378 vdd.n451 vdd.n450 0.0115
R1379 vdd.n508 vdd.n507 0.0113533
R1380 vdd.n624 vdd.n64 0.0113533
R1381 vdd.n468 vdd.n375 0.01106
R1382 vdd.n702 vdd.n34 0.01106
R1383 vdd.n483 vdd.n482 0.0109133
R1384 vdd.n600 vdd.n599 0.01062
R1385 vdd.n413 vdd.n412 0.0104733
R1386 vdd.n773 vdd.n12 0.0104733
R1387 vdd.n715 vdd.n714 0.0103267
R1388 vdd.n290 vdd 0.0102778
R1389 vdd.n515 vdd.n514 0.01018
R1390 vdd.n635 vdd.n62 0.01018
R1391 vdd.n479 vdd.n373 0.00988667
R1392 vdd.n677 vdd.n37 0.00988667
R1393 vdd.n680 vdd.n679 0.00974
R1394 vdd.n578 vdd.n577 0.00944667
R1395 vdd.n184 vdd.n183 0.00921287
R1396 vdd.n321 vdd.n184 0.00921287
R1397 vdd.n321 vdd.n320 0.00921287
R1398 vdd.n320 vdd.n318 0.00921287
R1399 vdd.n318 vdd.n185 0.00921287
R1400 vdd.n272 vdd.n185 0.00921287
R1401 vdd.n275 vdd.n272 0.00921287
R1402 vdd.n276 vdd.n275 0.00921287
R1403 vdd.n276 vdd.n270 0.00921287
R1404 vdd.n283 vdd.n270 0.00921287
R1405 vdd.n284 vdd.n283 0.00921287
R1406 vdd.n303 vdd.n284 0.00921287
R1407 vdd.n303 vdd.n302 0.00921287
R1408 vdd.n302 vdd.n298 0.00921287
R1409 vdd.n298 vdd.n297 0.00921287
R1410 vdd.n297 vdd.n285 0.00921287
R1411 vdd.n287 vdd.n285 0.00921287
R1412 vdd.n289 vdd.n287 0.00921287
R1413 vdd.n463 vdd.n384 0.00915333
R1414 vdd.n523 vdd.n522 0.00900667
R1415 vdd.n657 vdd.n656 0.00900667
R1416 vdd.n537 vdd.n536 0.00871333
R1417 vdd.n671 vdd.n670 0.00871333
R1418 vdd.n472 vdd.n471 0.00856667
R1419 vdd.n611 vdd.n610 0.00827333
R1420 vdd.n699 vdd.n698 0.00798
R1421 vdd.n664 vdd.n663 0.00783333
R1422 vdd.n664 vdd.n1 0.00783333
R1423 vdd.n558 vdd.n557 0.00783333
R1424 vdd.n558 vdd.n48 0.00783333
R1425 vdd.n531 vdd.n530 0.00783333
R1426 vdd.n650 vdd.n649 0.00783333
R1427 vdd.n530 vdd.n529 0.00754
R1428 vdd.n651 vdd.n650 0.00754
R1429 vdd.n698 vdd.n697 0.00739333
R1430 vdd.n610 vdd.n609 0.0071
R1431 vdd.n555 vdd.n355 0.00696745
R1432 vdd.n548 vdd.n354 0.00696745
R1433 vdd.n544 vdd.n353 0.00696745
R1434 vdd.n540 vdd.n352 0.00696745
R1435 vdd.n561 vdd.n49 0.00696745
R1436 vdd.n565 vdd.n50 0.00696745
R1437 vdd.n616 vdd.n51 0.00696745
R1438 vdd.n620 vdd.n52 0.00696745
R1439 vdd.n666 vdd.n6 0.00696745
R1440 vdd.n706 vdd.n5 0.00696745
R1441 vdd.n708 vdd.n4 0.00696745
R1442 vdd.n754 vdd.n3 0.00696745
R1443 vdd.n555 vdd.n554 0.00696745
R1444 vdd.n550 vdd.n354 0.00696745
R1445 vdd.n547 vdd.n353 0.00696745
R1446 vdd.n543 vdd.n352 0.00696745
R1447 vdd.n564 vdd.n49 0.00696745
R1448 vdd.n615 vdd.n50 0.00696745
R1449 vdd.n619 vdd.n51 0.00696745
R1450 vdd.n53 vdd.n52 0.00696745
R1451 vdd.n705 vdd.n6 0.00696745
R1452 vdd.n709 vdd.n5 0.00696745
R1453 vdd.n753 vdd.n4 0.00696745
R1454 vdd.n756 vdd.n3 0.00696745
R1455 vdd.n356 vdd.n90 0.00695265
R1456 vdd.n473 vdd.n472 0.00680667
R1457 vdd.n537 vdd.n367 0.00666
R1458 vdd.n670 vdd.n42 0.00666
R1459 vdd.n522 vdd.n520 0.00636667
R1460 vdd.n657 vdd.n56 0.00636667
R1461 vdd.n459 vdd.n384 0.00622
R1462 vdd.n779 vdd.n9 0.00607333
R1463 vdd.n176 vdd.n159 0.00606962
R1464 vdd.n266 vdd.n212 0.00603377
R1465 vdd.n784 vdd.n783 0.006
R1466 vdd.n577 vdd.n576 0.00592667
R1467 vdd.n679 vdd.n678 0.00563333
R1468 vdd.n476 vdd.n373 0.00548667
R1469 vdd.n681 vdd.n37 0.00548667
R1470 vdd.n114 vdd.n113 0.00538889
R1471 vdd.n114 vdd.n112 0.00538889
R1472 vdd.n117 vdd.n112 0.00538889
R1473 vdd.n118 vdd.n117 0.00538889
R1474 vdd.n119 vdd.n118 0.00538889
R1475 vdd.n120 vdd.n119 0.00538889
R1476 vdd.n121 vdd.n120 0.00538889
R1477 vdd.n121 vdd.n101 0.00538889
R1478 vdd.n124 vdd.n101 0.00538889
R1479 vdd.n124 vdd.n123 0.00538889
R1480 vdd.n123 vdd.n109 0.00538889
R1481 vdd.n338 vdd.n109 0.00538889
R1482 vdd.n338 vdd.n337 0.00538889
R1483 vdd.n337 vdd.n110 0.00538889
R1484 vdd.n334 vdd.n110 0.00538889
R1485 vdd.n334 vdd.n333 0.00538889
R1486 vdd.n333 vdd.n128 0.00538889
R1487 vdd.n164 vdd.n128 0.00538889
R1488 vdd.n165 vdd.n164 0.00538889
R1489 vdd.n166 vdd.n165 0.00538889
R1490 vdd.n167 vdd.n166 0.00538889
R1491 vdd.n167 vdd.n162 0.00538889
R1492 vdd.n170 vdd.n162 0.00538889
R1493 vdd.n171 vdd.n170 0.00538889
R1494 vdd.n172 vdd.n171 0.00538889
R1495 vdd.n173 vdd.n172 0.00538889
R1496 vdd.n174 vdd.n173 0.00538889
R1497 vdd.n174 vdd.n160 0.00538889
R1498 vdd.n177 vdd.n160 0.00538889
R1499 vdd.n178 vdd.n177 0.00538889
R1500 vdd.n182 vdd.n178 0.00538889
R1501 vdd.n182 vdd.n181 0.00538889
R1502 vdd.n181 vdd.n157 0.00538889
R1503 vdd.n323 vdd.n157 0.00538889
R1504 vdd.n323 vdd.n322 0.00538889
R1505 vdd.n322 vdd.n158 0.00538889
R1506 vdd.n319 vdd.n158 0.00538889
R1507 vdd.n319 vdd.n145 0.00538889
R1508 vdd.n317 vdd.n145 0.00538889
R1509 vdd.n317 vdd.n316 0.00538889
R1510 vdd.n316 vdd.n315 0.00538889
R1511 vdd.n315 vdd.n314 0.00538889
R1512 vdd.n314 vdd.n186 0.00538889
R1513 vdd.n273 vdd.n186 0.00538889
R1514 vdd.n274 vdd.n273 0.00538889
R1515 vdd.n274 vdd.n271 0.00538889
R1516 vdd.n277 vdd.n271 0.00538889
R1517 vdd.n278 vdd.n277 0.00538889
R1518 vdd.n279 vdd.n278 0.00538889
R1519 vdd.n280 vdd.n279 0.00538889
R1520 vdd.n282 vdd.n280 0.00538889
R1521 vdd.n282 vdd.n281 0.00538889
R1522 vdd.n281 vdd.n210 0.00538889
R1523 vdd.n305 vdd.n210 0.00538889
R1524 vdd.n305 vdd.n304 0.00538889
R1525 vdd.n304 vdd.n211 0.00538889
R1526 vdd.n301 vdd.n211 0.00538889
R1527 vdd.n301 vdd.n300 0.00538889
R1528 vdd.n300 vdd.n299 0.00538889
R1529 vdd.n299 vdd.n202 0.00538889
R1530 vdd.n296 vdd.n202 0.00538889
R1531 vdd.n296 vdd.n295 0.00538889
R1532 vdd.n295 vdd.n294 0.00538889
R1533 vdd.n294 vdd.n293 0.00538889
R1534 vdd.n293 vdd.n286 0.00538889
R1535 vdd.n291 vdd.n286 0.00538889
R1536 vdd.n291 vdd.n290 0.00538889
R1537 vdd.n514 vdd.n513 0.00519333
R1538 vdd.n632 vdd.n62 0.00519333
R1539 vdd.n716 vdd.n715 0.00504667
R1540 vdd.n412 vdd.n403 0.0049
R1541 vdd.n770 vdd.n12 0.0049
R1542 vdd.n183 vdd.n159 0.00485644
R1543 vdd.n289 vdd.n288 0.00485644
R1544 vdd.n288 vdd 0.00485644
R1545 vdd.n599 vdd.n598 0.00475333
R1546 vdd.n484 vdd.n483 0.00446
R1547 vdd.n469 vdd.n468 0.00431333
R1548 vdd.n702 vdd.n701 0.00431333
R1549 vdd.n414 vdd.n407 0.00416667
R1550 vdd.n783 vdd 0.00416667
R1551 vdd.n507 vdd.n506 0.00402
R1552 vdd.n625 vdd.n624 0.00402
R1553 vdd.n450 vdd.n449 0.00387333
R1554 vdd.n422 vdd.n401 0.00372667
R1555 vdd.n760 vdd.n759 0.00372667
R1556 vdd.n662 vdd.n48 0.00358
R1557 vdd.n504 vdd.n503 0.00358
R1558 vdd.n663 vdd.n662 0.00354333
R1559 vdd.n647 vdd.n646 0.00328667
R1560 vdd.n462 vdd.n461 0.00314
R1561 vdd.n694 vdd.n693 0.00314
R1562 vdd.n767 vdd.n766 0.00299333
R1563 vdd.n568 vdd.n82 0.00284667
R1564 vdd.n590 vdd.n71 0.00284667
R1565 vdd.n727 vdd.n22 0.0027
R1566 vdd.n429 vdd.n428 0.00255333
R1567 vdd.n744 vdd.n743 0.00255333
R1568 vdd.n339 vdd.n92 0.0025
R1569 vdd.n332 vdd.n92 0.0025
R1570 vdd.n332 vdd.n129 0.0025
R1571 vdd.n136 vdd.n129 0.0025
R1572 vdd.n326 vdd.n146 0.0025
R1573 vdd.n313 vdd.n146 0.0025
R1574 vdd.n313 vdd.n187 0.0025
R1575 vdd.n307 vdd.n194 0.0025
R1576 vdd.n310 vdd.n196 0.0025
R1577 vdd.n310 vdd.n203 0.0025
R1578 vdd.n292 vdd.n203 0.0025
R1579 vdd.n629 vdd.n628 0.00240667
R1580 vdd.n527 vdd.n526 0.00211333
R1581 vdd.n105 vdd.n96 0.00199909
R1582 vdd.n342 vdd.n105 0.00199909
R1583 vdd.n344 vdd.n97 0.00199909
R1584 vdd.n341 vdd.n97 0.00199909
R1585 vdd.n350 vdd.n98 0.00199909
R1586 vdd.n350 vdd.n102 0.00199909
R1587 vdd.n339 vdd.n108 0.00199909
R1588 vdd.n149 vdd.n136 0.00199909
R1589 vdd.n140 vdd.n135 0.00199909
R1590 vdd.n148 vdd.n140 0.00199909
R1591 vdd.n139 vdd.n134 0.00199909
R1592 vdd.n147 vdd.n139 0.00199909
R1593 vdd.n180 vdd.n133 0.00199909
R1594 vdd.n180 vdd.n138 0.00199909
R1595 vdd.n153 vdd.n132 0.00199909
R1596 vdd.n153 vdd.n144 0.00199909
R1597 vdd.n206 vdd.n191 0.00199909
R1598 vdd.n200 vdd.n191 0.00199909
R1599 vdd.n205 vdd.n190 0.00199909
R1600 vdd.n199 vdd.n190 0.00199909
R1601 vdd.n307 vdd.n209 0.00199909
R1602 vdd.n195 vdd.n194 0.00199909
R1603 vdd.n149 vdd.n141 0.00199909
R1604 vdd.n148 vdd.n142 0.00199909
R1605 vdd.n147 vdd.n143 0.00199909
R1606 vdd.n324 vdd.n138 0.00199909
R1607 vdd.n141 vdd.n135 0.00199909
R1608 vdd.n142 vdd.n134 0.00199909
R1609 vdd.n143 vdd.n133 0.00199909
R1610 vdd.n324 vdd.n132 0.00199909
R1611 vdd.n326 vdd.n144 0.00199909
R1612 vdd.n344 vdd.n95 0.00199909
R1613 vdd.n98 vdd.n94 0.00199909
R1614 vdd.n342 vdd.n95 0.00199909
R1615 vdd.n341 vdd.n94 0.00199909
R1616 vdd.n102 vdd.n93 0.00199909
R1617 vdd.n108 vdd.n93 0.00199909
R1618 vdd.n347 vdd.n96 0.00199909
R1619 vdd.n206 vdd.n187 0.00199909
R1620 vdd.n205 vdd.n192 0.00199909
R1621 vdd.n200 vdd.n192 0.00199909
R1622 vdd.n199 vdd.n193 0.00199909
R1623 vdd.n209 vdd.n193 0.00199909
R1624 vdd.n196 vdd.n195 0.00199909
R1625 vdd.n312 vdd.n130 0.00196667
R1626 vdd.n331 vdd.n330 0.00196667
R1627 vdd.n455 vdd.n454 0.00196667
R1628 vdd.n712 vdd.n25 0.00196667
R1629 vdd.n330 vdd.n329 0.00184933
R1630 vdd.n329 vdd.n130 0.001842
R1631 vdd.n424 vdd.n400 0.00182
R1632 vdd.n579 vdd.n77 0.00167333
R1633 vdd.n606 vdd.n588 0.00167333
R1634 vdd.n179 vdd.n151 0.00159978
R1635 vdd.n156 vdd.n155 0.00159978
R1636 vdd.n329 vdd.n131 0.00159978
R1637 vdd.n328 vdd.n327 0.00159978
R1638 vdd.n150 vdd.n137 0.00159978
R1639 vdd.n325 vdd.n152 0.00159978
R1640 vdd.n152 vdd.n150 0.00159978
R1641 vdd.n327 vdd.n137 0.00159978
R1642 vdd.n329 vdd.n328 0.00159978
R1643 vdd.n156 vdd.n131 0.00159978
R1644 vdd.n155 vdd.n151 0.00159978
R1645 vdd.n179 vdd.n154 0.00159978
R1646 vdd.n348 vdd.n99 0.00159978
R1647 vdd.n104 vdd.n100 0.00159978
R1648 vdd.n107 vdd.n100 0.00159978
R1649 vdd.n343 vdd.n340 0.00159978
R1650 vdd.n346 vdd.n343 0.00159978
R1651 vdd.n351 vdd.n91 0.00159978
R1652 vdd.n346 vdd.n345 0.00159978
R1653 vdd.n345 vdd.n91 0.00159978
R1654 vdd.n107 vdd.n103 0.00159978
R1655 vdd.n340 vdd.n103 0.00159978
R1656 vdd.n349 vdd.n348 0.00159978
R1657 vdd.n349 vdd.n104 0.00159978
R1658 vdd.n309 vdd.n208 0.00159978
R1659 vdd.n308 vdd.n198 0.00159978
R1660 vdd.n311 vdd.n188 0.00159978
R1661 vdd.n201 vdd.n189 0.00159978
R1662 vdd.n207 vdd.n204 0.00159978
R1663 vdd.n306 vdd.n0 0.00159978
R1664 vdd.n306 vdd.n207 0.00159978
R1665 vdd.n204 vdd.n201 0.00159978
R1666 vdd.n311 vdd.n189 0.00159978
R1667 vdd.n198 vdd.n188 0.00159978
R1668 vdd.n309 vdd.n308 0.00159978
R1669 vdd.n208 vdd.n197 0.00159978
R1670 vdd.n437 vdd.n436 0.00152667
R1671 vdd.n325 vdd 0.00140016
R1672 vdd.n662 vdd 0.00140016
R1673 vdd vdd.n351 0.00140016
R1674 vdd.n556 vdd 0.00140016
R1675 vdd vdd.n0 0.00140016
R1676 vdd.n784 vdd 0.00140016
R1677 vdd.n440 vdd.n439 0.00138
R1678 vdd.n750 vdd.n20 0.00138
R1679 vdd.n312 vdd.n311 0.001358
R1680 vdd.n331 vdd.n103 0.001358
R1681 vdd.n497 vdd.n492 0.00123333
R1682 vdd.n784 vdd.n1 0.00112333
R1683 vdd.n557 vdd.n556 0.00112333
R1684 vdd.n640 vdd.n639 0.00094
R1685 vdd.n447 vdd.n446 0.000793333
R1686 vdd.n720 vdd.n23 0.000793333
R1687 vdd.n739 vdd.n734 0.000646667
R1688 iovss.n87 iovss.n85 0.826084
R1689 iovss.n186 iovss.n1 0.826084
R1690 iovss.n86 iovss.n81 0.818682
R1691 iovss.n95 iovss.n80 0.818682
R1692 iovss.n96 iovss.n79 0.818682
R1693 iovss.n78 iovss.n74 0.818682
R1694 iovss.n103 iovss.n73 0.818682
R1695 iovss.n104 iovss.n72 0.818682
R1696 iovss.n71 iovss.n67 0.818682
R1697 iovss.n111 iovss.n66 0.818682
R1698 iovss.n112 iovss.n65 0.818682
R1699 iovss.n64 iovss.n60 0.818682
R1700 iovss.n119 iovss.n59 0.818682
R1701 iovss.n120 iovss.n58 0.818682
R1702 iovss.n57 iovss.n53 0.818682
R1703 iovss.n127 iovss.n52 0.818682
R1704 iovss.n128 iovss.n51 0.818682
R1705 iovss.n50 iovss.n46 0.818682
R1706 iovss.n135 iovss.n45 0.818682
R1707 iovss.n136 iovss.n44 0.818682
R1708 iovss.n43 iovss.n39 0.818682
R1709 iovss.n143 iovss.n38 0.818682
R1710 iovss.n144 iovss.n37 0.818682
R1711 iovss.n36 iovss.n32 0.818682
R1712 iovss.n151 iovss.n31 0.818682
R1713 iovss.n152 iovss.n30 0.818682
R1714 iovss.n29 iovss.n25 0.818682
R1715 iovss.n159 iovss.n24 0.818682
R1716 iovss.n160 iovss.n23 0.818682
R1717 iovss.n22 iovss.n18 0.818682
R1718 iovss.n167 iovss.n17 0.818682
R1719 iovss.n168 iovss.n16 0.818682
R1720 iovss.n15 iovss.n11 0.818682
R1721 iovss.n175 iovss.n10 0.818682
R1722 iovss.n176 iovss.n9 0.818682
R1723 iovss.n8 iovss.n4 0.818682
R1724 iovss.n183 iovss.n3 0.818682
R1725 iovss.n185 iovss.n184 0.818682
R1726 iovss.n183 iovss.n182 0.818682
R1727 iovss.n5 iovss.n4 0.818682
R1728 iovss.n177 iovss.n176 0.818682
R1729 iovss.n175 iovss.n174 0.818682
R1730 iovss.n12 iovss.n11 0.818682
R1731 iovss.n169 iovss.n168 0.818682
R1732 iovss.n167 iovss.n166 0.818682
R1733 iovss.n19 iovss.n18 0.818682
R1734 iovss.n161 iovss.n160 0.818682
R1735 iovss.n159 iovss.n158 0.818682
R1736 iovss.n26 iovss.n25 0.818682
R1737 iovss.n153 iovss.n152 0.818682
R1738 iovss.n151 iovss.n150 0.818682
R1739 iovss.n33 iovss.n32 0.818682
R1740 iovss.n145 iovss.n144 0.818682
R1741 iovss.n143 iovss.n142 0.818682
R1742 iovss.n40 iovss.n39 0.818682
R1743 iovss.n137 iovss.n136 0.818682
R1744 iovss.n135 iovss.n134 0.818682
R1745 iovss.n47 iovss.n46 0.818682
R1746 iovss.n129 iovss.n128 0.818682
R1747 iovss.n127 iovss.n126 0.818682
R1748 iovss.n54 iovss.n53 0.818682
R1749 iovss.n121 iovss.n120 0.818682
R1750 iovss.n119 iovss.n118 0.818682
R1751 iovss.n61 iovss.n60 0.818682
R1752 iovss.n113 iovss.n112 0.818682
R1753 iovss.n111 iovss.n110 0.818682
R1754 iovss.n68 iovss.n67 0.818682
R1755 iovss.n105 iovss.n104 0.818682
R1756 iovss.n103 iovss.n102 0.818682
R1757 iovss.n75 iovss.n74 0.818682
R1758 iovss.n97 iovss.n96 0.818682
R1759 iovss.n95 iovss.n94 0.818682
R1760 iovss.n82 iovss.n81 0.818682
R1761 iovss.n89 iovss.n88 0.818682
R1762 iovss.n3 iovss.n1 0.416993
R1763 iovss.n87 iovss.n86 0.416993
R1764 iovss.n85 iovss.n84 0.2005
R1765 iovss.n91 iovss.n90 0.2005
R1766 iovss.n93 iovss.n92 0.2005
R1767 iovss.n77 iovss.n76 0.2005
R1768 iovss.n99 iovss.n98 0.2005
R1769 iovss.n101 iovss.n100 0.2005
R1770 iovss.n70 iovss.n69 0.2005
R1771 iovss.n107 iovss.n106 0.2005
R1772 iovss.n109 iovss.n108 0.2005
R1773 iovss.n63 iovss.n62 0.2005
R1774 iovss.n115 iovss.n114 0.2005
R1775 iovss.n117 iovss.n116 0.2005
R1776 iovss.n56 iovss.n55 0.2005
R1777 iovss.n123 iovss.n122 0.2005
R1778 iovss.n125 iovss.n124 0.2005
R1779 iovss.n49 iovss.n48 0.2005
R1780 iovss.n131 iovss.n130 0.2005
R1781 iovss.n133 iovss.n132 0.2005
R1782 iovss.n42 iovss.n41 0.2005
R1783 iovss.n139 iovss.n138 0.2005
R1784 iovss.n141 iovss.n140 0.2005
R1785 iovss.n35 iovss.n34 0.2005
R1786 iovss.n147 iovss.n146 0.2005
R1787 iovss.n149 iovss.n148 0.2005
R1788 iovss.n28 iovss.n27 0.2005
R1789 iovss.n155 iovss.n154 0.2005
R1790 iovss.n157 iovss.n156 0.2005
R1791 iovss.n21 iovss.n20 0.2005
R1792 iovss.n163 iovss.n162 0.2005
R1793 iovss.n165 iovss.n164 0.2005
R1794 iovss.n14 iovss.n13 0.2005
R1795 iovss.n171 iovss.n170 0.2005
R1796 iovss.n173 iovss.n172 0.2005
R1797 iovss.n7 iovss.n6 0.2005
R1798 iovss.n179 iovss.n178 0.2005
R1799 iovss.n181 iovss.n180 0.2005
R1800 iovss.n2 iovss.n0 0.2005
R1801 iovss.n187 iovss.n186 0.2005
R1802 iovss iovss.n187 0.0778508
R1803 iovss.n83 iovss 0.0724109
R1804 iovss.n83 iovss 0.00862677
R1805 iovss.n84 iovss.n83 0.00808703
R1806 iovss.n8 iovss.n3 0.00740196
R1807 iovss.n9 iovss.n8 0.00740196
R1808 iovss.n10 iovss.n9 0.00740196
R1809 iovss.n15 iovss.n10 0.00740196
R1810 iovss.n16 iovss.n15 0.00740196
R1811 iovss.n17 iovss.n16 0.00740196
R1812 iovss.n22 iovss.n17 0.00740196
R1813 iovss.n23 iovss.n22 0.00740196
R1814 iovss.n24 iovss.n23 0.00740196
R1815 iovss.n29 iovss.n24 0.00740196
R1816 iovss.n30 iovss.n29 0.00740196
R1817 iovss.n31 iovss.n30 0.00740196
R1818 iovss.n36 iovss.n31 0.00740196
R1819 iovss.n37 iovss.n36 0.00740196
R1820 iovss.n38 iovss.n37 0.00740196
R1821 iovss.n43 iovss.n38 0.00740196
R1822 iovss.n44 iovss.n43 0.00740196
R1823 iovss.n45 iovss.n44 0.00740196
R1824 iovss.n50 iovss.n45 0.00740196
R1825 iovss.n51 iovss.n50 0.00740196
R1826 iovss.n52 iovss.n51 0.00740196
R1827 iovss.n57 iovss.n52 0.00740196
R1828 iovss.n58 iovss.n57 0.00740196
R1829 iovss.n59 iovss.n58 0.00740196
R1830 iovss.n64 iovss.n59 0.00740196
R1831 iovss.n65 iovss.n64 0.00740196
R1832 iovss.n66 iovss.n65 0.00740196
R1833 iovss.n71 iovss.n66 0.00740196
R1834 iovss.n72 iovss.n71 0.00740196
R1835 iovss.n73 iovss.n72 0.00740196
R1836 iovss.n78 iovss.n73 0.00740196
R1837 iovss.n79 iovss.n78 0.00740196
R1838 iovss.n80 iovss.n79 0.00740196
R1839 iovss.n86 iovss.n80 0.00740196
R1840 iovss.n184 iovss.n183 0.00740196
R1841 iovss.n183 iovss.n4 0.00740196
R1842 iovss.n176 iovss.n4 0.00740196
R1843 iovss.n176 iovss.n175 0.00740196
R1844 iovss.n175 iovss.n11 0.00740196
R1845 iovss.n168 iovss.n11 0.00740196
R1846 iovss.n168 iovss.n167 0.00740196
R1847 iovss.n167 iovss.n18 0.00740196
R1848 iovss.n160 iovss.n18 0.00740196
R1849 iovss.n160 iovss.n159 0.00740196
R1850 iovss.n159 iovss.n25 0.00740196
R1851 iovss.n152 iovss.n25 0.00740196
R1852 iovss.n152 iovss.n151 0.00740196
R1853 iovss.n151 iovss.n32 0.00740196
R1854 iovss.n144 iovss.n32 0.00740196
R1855 iovss.n144 iovss.n143 0.00740196
R1856 iovss.n143 iovss.n39 0.00740196
R1857 iovss.n136 iovss.n39 0.00740196
R1858 iovss.n136 iovss.n135 0.00740196
R1859 iovss.n135 iovss.n46 0.00740196
R1860 iovss.n128 iovss.n46 0.00740196
R1861 iovss.n128 iovss.n127 0.00740196
R1862 iovss.n127 iovss.n53 0.00740196
R1863 iovss.n120 iovss.n53 0.00740196
R1864 iovss.n120 iovss.n119 0.00740196
R1865 iovss.n119 iovss.n60 0.00740196
R1866 iovss.n112 iovss.n60 0.00740196
R1867 iovss.n112 iovss.n111 0.00740196
R1868 iovss.n111 iovss.n67 0.00740196
R1869 iovss.n104 iovss.n67 0.00740196
R1870 iovss.n104 iovss.n103 0.00740196
R1871 iovss.n103 iovss.n74 0.00740196
R1872 iovss.n96 iovss.n74 0.00740196
R1873 iovss.n96 iovss.n95 0.00740196
R1874 iovss.n95 iovss.n81 0.00740196
R1875 iovss.n88 iovss.n81 0.00740196
R1876 iovss.n88 iovss.n87 0.00442211
R1877 iovss.n184 iovss.n1 0.00442211
R1878 iovss.n186 iovss.n185 0.00395098
R1879 iovss.n185 iovss.n2 0.00395098
R1880 iovss.n182 iovss.n2 0.00395098
R1881 iovss.n182 iovss.n181 0.00395098
R1882 iovss.n181 iovss.n5 0.00395098
R1883 iovss.n178 iovss.n5 0.00395098
R1884 iovss.n178 iovss.n177 0.00395098
R1885 iovss.n177 iovss.n7 0.00395098
R1886 iovss.n174 iovss.n7 0.00395098
R1887 iovss.n174 iovss.n173 0.00395098
R1888 iovss.n173 iovss.n12 0.00395098
R1889 iovss.n170 iovss.n12 0.00395098
R1890 iovss.n170 iovss.n169 0.00395098
R1891 iovss.n169 iovss.n14 0.00395098
R1892 iovss.n166 iovss.n14 0.00395098
R1893 iovss.n166 iovss.n165 0.00395098
R1894 iovss.n165 iovss.n19 0.00395098
R1895 iovss.n162 iovss.n19 0.00395098
R1896 iovss.n162 iovss.n161 0.00395098
R1897 iovss.n161 iovss.n21 0.00395098
R1898 iovss.n158 iovss.n21 0.00395098
R1899 iovss.n158 iovss.n157 0.00395098
R1900 iovss.n157 iovss.n26 0.00395098
R1901 iovss.n154 iovss.n26 0.00395098
R1902 iovss.n154 iovss.n153 0.00395098
R1903 iovss.n153 iovss.n28 0.00395098
R1904 iovss.n150 iovss.n28 0.00395098
R1905 iovss.n150 iovss.n149 0.00395098
R1906 iovss.n149 iovss.n33 0.00395098
R1907 iovss.n146 iovss.n33 0.00395098
R1908 iovss.n146 iovss.n145 0.00395098
R1909 iovss.n145 iovss.n35 0.00395098
R1910 iovss.n142 iovss.n35 0.00395098
R1911 iovss.n142 iovss.n141 0.00395098
R1912 iovss.n141 iovss.n40 0.00395098
R1913 iovss.n138 iovss.n40 0.00395098
R1914 iovss.n138 iovss.n137 0.00395098
R1915 iovss.n137 iovss.n42 0.00395098
R1916 iovss.n134 iovss.n42 0.00395098
R1917 iovss.n134 iovss.n133 0.00395098
R1918 iovss.n133 iovss.n47 0.00395098
R1919 iovss.n130 iovss.n47 0.00395098
R1920 iovss.n130 iovss.n129 0.00395098
R1921 iovss.n129 iovss.n49 0.00395098
R1922 iovss.n126 iovss.n49 0.00395098
R1923 iovss.n126 iovss.n125 0.00395098
R1924 iovss.n125 iovss.n54 0.00395098
R1925 iovss.n122 iovss.n54 0.00395098
R1926 iovss.n122 iovss.n121 0.00395098
R1927 iovss.n121 iovss.n56 0.00395098
R1928 iovss.n118 iovss.n56 0.00395098
R1929 iovss.n118 iovss.n117 0.00395098
R1930 iovss.n117 iovss.n61 0.00395098
R1931 iovss.n114 iovss.n61 0.00395098
R1932 iovss.n114 iovss.n113 0.00395098
R1933 iovss.n113 iovss.n63 0.00395098
R1934 iovss.n110 iovss.n63 0.00395098
R1935 iovss.n110 iovss.n109 0.00395098
R1936 iovss.n109 iovss.n68 0.00395098
R1937 iovss.n106 iovss.n68 0.00395098
R1938 iovss.n106 iovss.n105 0.00395098
R1939 iovss.n105 iovss.n70 0.00395098
R1940 iovss.n102 iovss.n70 0.00395098
R1941 iovss.n102 iovss.n101 0.00395098
R1942 iovss.n101 iovss.n75 0.00395098
R1943 iovss.n98 iovss.n75 0.00395098
R1944 iovss.n98 iovss.n97 0.00395098
R1945 iovss.n97 iovss.n77 0.00395098
R1946 iovss.n94 iovss.n77 0.00395098
R1947 iovss.n94 iovss.n93 0.00395098
R1948 iovss.n93 iovss.n82 0.00395098
R1949 iovss.n90 iovss.n82 0.00395098
R1950 iovss.n90 iovss.n89 0.00395098
R1951 iovss.n89 iovss.n85 0.00395098
R1952 iovss.n187 iovss.n0 0.00191176
R1953 iovss.n180 iovss.n0 0.00191176
R1954 iovss.n180 iovss.n179 0.00191176
R1955 iovss.n179 iovss.n6 0.00191176
R1956 iovss.n172 iovss.n6 0.00191176
R1957 iovss.n172 iovss.n171 0.00191176
R1958 iovss.n171 iovss.n13 0.00191176
R1959 iovss.n164 iovss.n13 0.00191176
R1960 iovss.n164 iovss.n163 0.00191176
R1961 iovss.n163 iovss.n20 0.00191176
R1962 iovss.n156 iovss.n20 0.00191176
R1963 iovss.n156 iovss.n155 0.00191176
R1964 iovss.n155 iovss.n27 0.00191176
R1965 iovss.n148 iovss.n27 0.00191176
R1966 iovss.n148 iovss.n147 0.00191176
R1967 iovss.n147 iovss.n34 0.00191176
R1968 iovss.n140 iovss.n34 0.00191176
R1969 iovss.n140 iovss.n139 0.00191176
R1970 iovss.n139 iovss.n41 0.00191176
R1971 iovss.n132 iovss.n41 0.00191176
R1972 iovss.n132 iovss.n131 0.00191176
R1973 iovss.n131 iovss.n48 0.00191176
R1974 iovss.n124 iovss.n48 0.00191176
R1975 iovss.n124 iovss.n123 0.00191176
R1976 iovss.n123 iovss.n55 0.00191176
R1977 iovss.n116 iovss.n55 0.00191176
R1978 iovss.n116 iovss.n115 0.00191176
R1979 iovss.n115 iovss.n62 0.00191176
R1980 iovss.n108 iovss.n62 0.00191176
R1981 iovss.n108 iovss.n107 0.00191176
R1982 iovss.n107 iovss.n69 0.00191176
R1983 iovss.n100 iovss.n69 0.00191176
R1984 iovss.n100 iovss.n99 0.00191176
R1985 iovss.n99 iovss.n76 0.00191176
R1986 iovss.n92 iovss.n76 0.00191176
R1987 iovss.n92 iovss.n91 0.00191176
R1988 iovss.n91 iovss.n84 0.00191176
R1989 sg13g2_RCClampInverter_0.in.n0 sg13g2_RCClampInverter_0.in.t1 10.5567
R1990 sg13g2_RCClampInverter_0.in.n0 sg13g2_RCClampInverter_0.in.t2 10.286
R1991 sg13g2_RCClampInverter_0.in.n1 sg13g2_RCClampInverter_0.in.t0 5.0005
R1992 sg13g2_RCClampInverter_0.in.n1 sg13g2_RCClampInverter_0.in 3.73153
R1993 sg13g2_RCClampInverter_0.in sg13g2_RCClampInverter_0.in.n1 0.0214524
R1994 sg13g2_RCClampInverter_0.in sg13g2_RCClampInverter_0.in.n0 0.00107971
R1995 iovdd.n87 iovdd.n85 0.826084
R1996 iovdd.n186 iovdd.n1 0.826084
R1997 iovdd.n86 iovdd.n81 0.818682
R1998 iovdd.n95 iovdd.n80 0.818682
R1999 iovdd.n96 iovdd.n79 0.818682
R2000 iovdd.n78 iovdd.n74 0.818682
R2001 iovdd.n103 iovdd.n73 0.818682
R2002 iovdd.n104 iovdd.n72 0.818682
R2003 iovdd.n71 iovdd.n67 0.818682
R2004 iovdd.n111 iovdd.n66 0.818682
R2005 iovdd.n112 iovdd.n65 0.818682
R2006 iovdd.n64 iovdd.n60 0.818682
R2007 iovdd.n119 iovdd.n59 0.818682
R2008 iovdd.n120 iovdd.n58 0.818682
R2009 iovdd.n57 iovdd.n53 0.818682
R2010 iovdd.n127 iovdd.n52 0.818682
R2011 iovdd.n128 iovdd.n51 0.818682
R2012 iovdd.n50 iovdd.n46 0.818682
R2013 iovdd.n135 iovdd.n45 0.818682
R2014 iovdd.n136 iovdd.n44 0.818682
R2015 iovdd.n43 iovdd.n39 0.818682
R2016 iovdd.n143 iovdd.n38 0.818682
R2017 iovdd.n144 iovdd.n37 0.818682
R2018 iovdd.n36 iovdd.n32 0.818682
R2019 iovdd.n151 iovdd.n31 0.818682
R2020 iovdd.n152 iovdd.n30 0.818682
R2021 iovdd.n29 iovdd.n25 0.818682
R2022 iovdd.n159 iovdd.n24 0.818682
R2023 iovdd.n160 iovdd.n23 0.818682
R2024 iovdd.n22 iovdd.n18 0.818682
R2025 iovdd.n167 iovdd.n17 0.818682
R2026 iovdd.n168 iovdd.n16 0.818682
R2027 iovdd.n15 iovdd.n11 0.818682
R2028 iovdd.n175 iovdd.n10 0.818682
R2029 iovdd.n176 iovdd.n9 0.818682
R2030 iovdd.n8 iovdd.n4 0.818682
R2031 iovdd.n183 iovdd.n3 0.818682
R2032 iovdd.n185 iovdd.n184 0.818682
R2033 iovdd.n183 iovdd.n182 0.818682
R2034 iovdd.n5 iovdd.n4 0.818682
R2035 iovdd.n177 iovdd.n176 0.818682
R2036 iovdd.n175 iovdd.n174 0.818682
R2037 iovdd.n12 iovdd.n11 0.818682
R2038 iovdd.n169 iovdd.n168 0.818682
R2039 iovdd.n167 iovdd.n166 0.818682
R2040 iovdd.n19 iovdd.n18 0.818682
R2041 iovdd.n161 iovdd.n160 0.818682
R2042 iovdd.n159 iovdd.n158 0.818682
R2043 iovdd.n26 iovdd.n25 0.818682
R2044 iovdd.n153 iovdd.n152 0.818682
R2045 iovdd.n151 iovdd.n150 0.818682
R2046 iovdd.n33 iovdd.n32 0.818682
R2047 iovdd.n145 iovdd.n144 0.818682
R2048 iovdd.n143 iovdd.n142 0.818682
R2049 iovdd.n40 iovdd.n39 0.818682
R2050 iovdd.n137 iovdd.n136 0.818682
R2051 iovdd.n135 iovdd.n134 0.818682
R2052 iovdd.n47 iovdd.n46 0.818682
R2053 iovdd.n129 iovdd.n128 0.818682
R2054 iovdd.n127 iovdd.n126 0.818682
R2055 iovdd.n54 iovdd.n53 0.818682
R2056 iovdd.n121 iovdd.n120 0.818682
R2057 iovdd.n119 iovdd.n118 0.818682
R2058 iovdd.n61 iovdd.n60 0.818682
R2059 iovdd.n113 iovdd.n112 0.818682
R2060 iovdd.n111 iovdd.n110 0.818682
R2061 iovdd.n68 iovdd.n67 0.818682
R2062 iovdd.n105 iovdd.n104 0.818682
R2063 iovdd.n103 iovdd.n102 0.818682
R2064 iovdd.n75 iovdd.n74 0.818682
R2065 iovdd.n97 iovdd.n96 0.818682
R2066 iovdd.n95 iovdd.n94 0.818682
R2067 iovdd.n82 iovdd.n81 0.818682
R2068 iovdd.n89 iovdd.n88 0.818682
R2069 iovdd.n3 iovdd.n1 0.416993
R2070 iovdd.n87 iovdd.n86 0.416993
R2071 iovdd.n85 iovdd.n84 0.2005
R2072 iovdd.n91 iovdd.n90 0.2005
R2073 iovdd.n93 iovdd.n92 0.2005
R2074 iovdd.n77 iovdd.n76 0.2005
R2075 iovdd.n99 iovdd.n98 0.2005
R2076 iovdd.n101 iovdd.n100 0.2005
R2077 iovdd.n70 iovdd.n69 0.2005
R2078 iovdd.n107 iovdd.n106 0.2005
R2079 iovdd.n109 iovdd.n108 0.2005
R2080 iovdd.n63 iovdd.n62 0.2005
R2081 iovdd.n115 iovdd.n114 0.2005
R2082 iovdd.n117 iovdd.n116 0.2005
R2083 iovdd.n56 iovdd.n55 0.2005
R2084 iovdd.n123 iovdd.n122 0.2005
R2085 iovdd.n125 iovdd.n124 0.2005
R2086 iovdd.n49 iovdd.n48 0.2005
R2087 iovdd.n131 iovdd.n130 0.2005
R2088 iovdd.n133 iovdd.n132 0.2005
R2089 iovdd.n42 iovdd.n41 0.2005
R2090 iovdd.n139 iovdd.n138 0.2005
R2091 iovdd.n141 iovdd.n140 0.2005
R2092 iovdd.n35 iovdd.n34 0.2005
R2093 iovdd.n147 iovdd.n146 0.2005
R2094 iovdd.n149 iovdd.n148 0.2005
R2095 iovdd.n28 iovdd.n27 0.2005
R2096 iovdd.n155 iovdd.n154 0.2005
R2097 iovdd.n157 iovdd.n156 0.2005
R2098 iovdd.n21 iovdd.n20 0.2005
R2099 iovdd.n163 iovdd.n162 0.2005
R2100 iovdd.n165 iovdd.n164 0.2005
R2101 iovdd.n14 iovdd.n13 0.2005
R2102 iovdd.n171 iovdd.n170 0.2005
R2103 iovdd.n173 iovdd.n172 0.2005
R2104 iovdd.n7 iovdd.n6 0.2005
R2105 iovdd.n179 iovdd.n178 0.2005
R2106 iovdd.n181 iovdd.n180 0.2005
R2107 iovdd.n2 iovdd.n0 0.2005
R2108 iovdd.n187 iovdd.n186 0.2005
R2109 iovdd iovdd.n187 0.0778508
R2110 iovdd.n83 iovdd 0.0724109
R2111 iovdd.n83 iovdd 0.00862677
R2112 iovdd.n84 iovdd.n83 0.00808703
R2113 iovdd.n8 iovdd.n3 0.00740196
R2114 iovdd.n9 iovdd.n8 0.00740196
R2115 iovdd.n10 iovdd.n9 0.00740196
R2116 iovdd.n15 iovdd.n10 0.00740196
R2117 iovdd.n16 iovdd.n15 0.00740196
R2118 iovdd.n17 iovdd.n16 0.00740196
R2119 iovdd.n22 iovdd.n17 0.00740196
R2120 iovdd.n23 iovdd.n22 0.00740196
R2121 iovdd.n24 iovdd.n23 0.00740196
R2122 iovdd.n29 iovdd.n24 0.00740196
R2123 iovdd.n30 iovdd.n29 0.00740196
R2124 iovdd.n31 iovdd.n30 0.00740196
R2125 iovdd.n36 iovdd.n31 0.00740196
R2126 iovdd.n37 iovdd.n36 0.00740196
R2127 iovdd.n38 iovdd.n37 0.00740196
R2128 iovdd.n43 iovdd.n38 0.00740196
R2129 iovdd.n44 iovdd.n43 0.00740196
R2130 iovdd.n45 iovdd.n44 0.00740196
R2131 iovdd.n50 iovdd.n45 0.00740196
R2132 iovdd.n51 iovdd.n50 0.00740196
R2133 iovdd.n52 iovdd.n51 0.00740196
R2134 iovdd.n57 iovdd.n52 0.00740196
R2135 iovdd.n58 iovdd.n57 0.00740196
R2136 iovdd.n59 iovdd.n58 0.00740196
R2137 iovdd.n64 iovdd.n59 0.00740196
R2138 iovdd.n65 iovdd.n64 0.00740196
R2139 iovdd.n66 iovdd.n65 0.00740196
R2140 iovdd.n71 iovdd.n66 0.00740196
R2141 iovdd.n72 iovdd.n71 0.00740196
R2142 iovdd.n73 iovdd.n72 0.00740196
R2143 iovdd.n78 iovdd.n73 0.00740196
R2144 iovdd.n79 iovdd.n78 0.00740196
R2145 iovdd.n80 iovdd.n79 0.00740196
R2146 iovdd.n86 iovdd.n80 0.00740196
R2147 iovdd.n184 iovdd.n183 0.00740196
R2148 iovdd.n183 iovdd.n4 0.00740196
R2149 iovdd.n176 iovdd.n4 0.00740196
R2150 iovdd.n176 iovdd.n175 0.00740196
R2151 iovdd.n175 iovdd.n11 0.00740196
R2152 iovdd.n168 iovdd.n11 0.00740196
R2153 iovdd.n168 iovdd.n167 0.00740196
R2154 iovdd.n167 iovdd.n18 0.00740196
R2155 iovdd.n160 iovdd.n18 0.00740196
R2156 iovdd.n160 iovdd.n159 0.00740196
R2157 iovdd.n159 iovdd.n25 0.00740196
R2158 iovdd.n152 iovdd.n25 0.00740196
R2159 iovdd.n152 iovdd.n151 0.00740196
R2160 iovdd.n151 iovdd.n32 0.00740196
R2161 iovdd.n144 iovdd.n32 0.00740196
R2162 iovdd.n144 iovdd.n143 0.00740196
R2163 iovdd.n143 iovdd.n39 0.00740196
R2164 iovdd.n136 iovdd.n39 0.00740196
R2165 iovdd.n136 iovdd.n135 0.00740196
R2166 iovdd.n135 iovdd.n46 0.00740196
R2167 iovdd.n128 iovdd.n46 0.00740196
R2168 iovdd.n128 iovdd.n127 0.00740196
R2169 iovdd.n127 iovdd.n53 0.00740196
R2170 iovdd.n120 iovdd.n53 0.00740196
R2171 iovdd.n120 iovdd.n119 0.00740196
R2172 iovdd.n119 iovdd.n60 0.00740196
R2173 iovdd.n112 iovdd.n60 0.00740196
R2174 iovdd.n112 iovdd.n111 0.00740196
R2175 iovdd.n111 iovdd.n67 0.00740196
R2176 iovdd.n104 iovdd.n67 0.00740196
R2177 iovdd.n104 iovdd.n103 0.00740196
R2178 iovdd.n103 iovdd.n74 0.00740196
R2179 iovdd.n96 iovdd.n74 0.00740196
R2180 iovdd.n96 iovdd.n95 0.00740196
R2181 iovdd.n95 iovdd.n81 0.00740196
R2182 iovdd.n88 iovdd.n81 0.00740196
R2183 iovdd.n88 iovdd.n87 0.00442211
R2184 iovdd.n184 iovdd.n1 0.00442211
R2185 iovdd.n186 iovdd.n185 0.00395098
R2186 iovdd.n185 iovdd.n2 0.00395098
R2187 iovdd.n182 iovdd.n2 0.00395098
R2188 iovdd.n182 iovdd.n181 0.00395098
R2189 iovdd.n181 iovdd.n5 0.00395098
R2190 iovdd.n178 iovdd.n5 0.00395098
R2191 iovdd.n178 iovdd.n177 0.00395098
R2192 iovdd.n177 iovdd.n7 0.00395098
R2193 iovdd.n174 iovdd.n7 0.00395098
R2194 iovdd.n174 iovdd.n173 0.00395098
R2195 iovdd.n173 iovdd.n12 0.00395098
R2196 iovdd.n170 iovdd.n12 0.00395098
R2197 iovdd.n170 iovdd.n169 0.00395098
R2198 iovdd.n169 iovdd.n14 0.00395098
R2199 iovdd.n166 iovdd.n14 0.00395098
R2200 iovdd.n166 iovdd.n165 0.00395098
R2201 iovdd.n165 iovdd.n19 0.00395098
R2202 iovdd.n162 iovdd.n19 0.00395098
R2203 iovdd.n162 iovdd.n161 0.00395098
R2204 iovdd.n161 iovdd.n21 0.00395098
R2205 iovdd.n158 iovdd.n21 0.00395098
R2206 iovdd.n158 iovdd.n157 0.00395098
R2207 iovdd.n157 iovdd.n26 0.00395098
R2208 iovdd.n154 iovdd.n26 0.00395098
R2209 iovdd.n154 iovdd.n153 0.00395098
R2210 iovdd.n153 iovdd.n28 0.00395098
R2211 iovdd.n150 iovdd.n28 0.00395098
R2212 iovdd.n150 iovdd.n149 0.00395098
R2213 iovdd.n149 iovdd.n33 0.00395098
R2214 iovdd.n146 iovdd.n33 0.00395098
R2215 iovdd.n146 iovdd.n145 0.00395098
R2216 iovdd.n145 iovdd.n35 0.00395098
R2217 iovdd.n142 iovdd.n35 0.00395098
R2218 iovdd.n142 iovdd.n141 0.00395098
R2219 iovdd.n141 iovdd.n40 0.00395098
R2220 iovdd.n138 iovdd.n40 0.00395098
R2221 iovdd.n138 iovdd.n137 0.00395098
R2222 iovdd.n137 iovdd.n42 0.00395098
R2223 iovdd.n134 iovdd.n42 0.00395098
R2224 iovdd.n134 iovdd.n133 0.00395098
R2225 iovdd.n133 iovdd.n47 0.00395098
R2226 iovdd.n130 iovdd.n47 0.00395098
R2227 iovdd.n130 iovdd.n129 0.00395098
R2228 iovdd.n129 iovdd.n49 0.00395098
R2229 iovdd.n126 iovdd.n49 0.00395098
R2230 iovdd.n126 iovdd.n125 0.00395098
R2231 iovdd.n125 iovdd.n54 0.00395098
R2232 iovdd.n122 iovdd.n54 0.00395098
R2233 iovdd.n122 iovdd.n121 0.00395098
R2234 iovdd.n121 iovdd.n56 0.00395098
R2235 iovdd.n118 iovdd.n56 0.00395098
R2236 iovdd.n118 iovdd.n117 0.00395098
R2237 iovdd.n117 iovdd.n61 0.00395098
R2238 iovdd.n114 iovdd.n61 0.00395098
R2239 iovdd.n114 iovdd.n113 0.00395098
R2240 iovdd.n113 iovdd.n63 0.00395098
R2241 iovdd.n110 iovdd.n63 0.00395098
R2242 iovdd.n110 iovdd.n109 0.00395098
R2243 iovdd.n109 iovdd.n68 0.00395098
R2244 iovdd.n106 iovdd.n68 0.00395098
R2245 iovdd.n106 iovdd.n105 0.00395098
R2246 iovdd.n105 iovdd.n70 0.00395098
R2247 iovdd.n102 iovdd.n70 0.00395098
R2248 iovdd.n102 iovdd.n101 0.00395098
R2249 iovdd.n101 iovdd.n75 0.00395098
R2250 iovdd.n98 iovdd.n75 0.00395098
R2251 iovdd.n98 iovdd.n97 0.00395098
R2252 iovdd.n97 iovdd.n77 0.00395098
R2253 iovdd.n94 iovdd.n77 0.00395098
R2254 iovdd.n94 iovdd.n93 0.00395098
R2255 iovdd.n93 iovdd.n82 0.00395098
R2256 iovdd.n90 iovdd.n82 0.00395098
R2257 iovdd.n90 iovdd.n89 0.00395098
R2258 iovdd.n89 iovdd.n85 0.00395098
R2259 iovdd.n187 iovdd.n0 0.00191176
R2260 iovdd.n180 iovdd.n0 0.00191176
R2261 iovdd.n180 iovdd.n179 0.00191176
R2262 iovdd.n179 iovdd.n6 0.00191176
R2263 iovdd.n172 iovdd.n6 0.00191176
R2264 iovdd.n172 iovdd.n171 0.00191176
R2265 iovdd.n171 iovdd.n13 0.00191176
R2266 iovdd.n164 iovdd.n13 0.00191176
R2267 iovdd.n164 iovdd.n163 0.00191176
R2268 iovdd.n163 iovdd.n20 0.00191176
R2269 iovdd.n156 iovdd.n20 0.00191176
R2270 iovdd.n156 iovdd.n155 0.00191176
R2271 iovdd.n155 iovdd.n27 0.00191176
R2272 iovdd.n148 iovdd.n27 0.00191176
R2273 iovdd.n148 iovdd.n147 0.00191176
R2274 iovdd.n147 iovdd.n34 0.00191176
R2275 iovdd.n140 iovdd.n34 0.00191176
R2276 iovdd.n140 iovdd.n139 0.00191176
R2277 iovdd.n139 iovdd.n41 0.00191176
R2278 iovdd.n132 iovdd.n41 0.00191176
R2279 iovdd.n132 iovdd.n131 0.00191176
R2280 iovdd.n131 iovdd.n48 0.00191176
R2281 iovdd.n124 iovdd.n48 0.00191176
R2282 iovdd.n124 iovdd.n123 0.00191176
R2283 iovdd.n123 iovdd.n55 0.00191176
R2284 iovdd.n116 iovdd.n55 0.00191176
R2285 iovdd.n116 iovdd.n115 0.00191176
R2286 iovdd.n115 iovdd.n62 0.00191176
R2287 iovdd.n108 iovdd.n62 0.00191176
R2288 iovdd.n108 iovdd.n107 0.00191176
R2289 iovdd.n107 iovdd.n69 0.00191176
R2290 iovdd.n100 iovdd.n69 0.00191176
R2291 iovdd.n100 iovdd.n99 0.00191176
R2292 iovdd.n99 iovdd.n76 0.00191176
R2293 iovdd.n92 iovdd.n76 0.00191176
R2294 iovdd.n92 iovdd.n91 0.00191176
R2295 iovdd.n91 iovdd.n84 0.00191176
C0 a_6085_7542# a_6415_7542# 0.37213f
C1 a_5755_7542# a_5425_7542# 0.37213f
C2 a_4765_7542# a_4435_7542# 0.37213f
C3 a_6745_7542# a_7075_7542# 0.37213f
C4 a_10705_7542# a_10375_7542# 0.37213f
C5 a_11695_7542# a_12025_7542# 0.37213f
C6 a_3775_7542# a_4105_7542# 0.37213f
C7 vdd w_n124_1076# 6.51124f
C8 a_9055_7542# a_9385_7542# 0.37213f
C9 sg13g2_RCClampInverter_0.out w_n124_1076# 2.16343f
C10 sg13g2_RCClampInverter_0.out vdd 89.81529f
C11 a_7405_7542# a_7735_7542# 0.37213f
C12 sg13g2_RCClampInverter_0.in w_n124_1076# 3.24089f
C13 sg13g2_RCClampInverter_0.in vdd 31.5477f
C14 iovdd w_n124_1076# 1.22195f
C15 vdd iovdd 0.12505p
C16 sg13g2_RCClampInverter_0.in sg13g2_RCClampInverter_0.out 21.6731f
C17 sg13g2_RCClampInverter_0.out iovdd 43.9772f
C18 a_4105_7542# a_4435_7542# 0.37213f
C19 a_10045_7542# a_10375_7542# 0.37213f
C20 a_6745_7542# a_6415_7542# 0.37213f
C21 a_9715_7542# a_10045_7542# 0.37213f
C22 sg13g2_RCClampInverter_0.in iovdd 55.64351f
C23 a_9715_7542# a_9385_7542# 0.37213f
C24 a_4765_7542# a_5095_7542# 0.37213f
C25 a_10705_7542# a_11035_7542# 0.37213f
C26 a_11695_7542# a_11365_7542# 0.37213f
C27 a_8725_7542# a_9055_7542# 0.37213f
C28 a_8395_7542# a_8725_7542# 0.37213f
C29 a_8065_7542# a_8395_7542# 0.37213f
C30 a_11365_7542# a_11035_7542# 0.37213f
C31 a_7405_7542# a_7075_7542# 0.37213f
C32 a_5095_7542# a_5425_7542# 0.37213f
C33 a_8065_7542# a_7735_7542# 0.37213f
C34 a_6085_7542# a_5755_7542# 0.37213f
C35 iovdd iovss 67.28207f
C36 vdd iovss 0.69054p
C37 a_12025_7542# iovss 3.53966f $ **FLOATING
C38 a_11695_7456# iovss 0.45487f
C39 a_11695_7542# iovss 3.04229f $ **FLOATING
C40 a_11365_7542# iovss 3.04218f $ **FLOATING
C41 a_11365_11542# iovss 0.41716f
C42 a_11035_7456# iovss 0.43382f
C43 a_11035_7542# iovss 3.04229f $ **FLOATING
C44 a_10705_7542# iovss 3.04218f $ **FLOATING
C45 a_10705_11542# iovss 0.41716f
C46 a_10375_7456# iovss 0.43383f
C47 a_10375_7542# iovss 3.04226f $ **FLOATING
C48 a_10045_7542# iovss 3.04218f $ **FLOATING
C49 a_10045_11542# iovss 0.41716f
C50 a_9715_7456# iovss 0.43386f
C51 a_9715_7542# iovss 3.04218f $ **FLOATING
C52 a_9385_7542# iovss 3.04218f $ **FLOATING
C53 a_9385_11542# iovss 0.41716f
C54 a_9055_7456# iovss 0.43385f
C55 a_9055_7542# iovss 3.04218f $ **FLOATING
C56 a_8725_7542# iovss 3.04229f $ **FLOATING
C57 a_8725_11542# iovss 0.41716f
C58 a_8395_7456# iovss 0.43382f
C59 a_8395_7542# iovss 3.04218f $ **FLOATING
C60 a_8065_7542# iovss 3.04229f $ **FLOATING
C61 a_8065_11542# iovss 0.41716f
C62 a_7735_7456# iovss 0.43382f
C63 a_7735_7542# iovss 3.04218f $ **FLOATING
C64 a_7405_7542# iovss 3.04229f $ **FLOATING
C65 a_7405_11542# iovss 0.41716f
C66 a_7075_7456# iovss 0.43384f
C67 a_7075_7542# iovss 3.04218f $ **FLOATING
C68 a_6745_7542# iovss 3.04224f $ **FLOATING
C69 a_6745_11542# iovss 0.41716f
C70 a_6415_7456# iovss 0.43388f
C71 a_6415_7542# iovss 3.04218f $ **FLOATING
C72 a_6085_7542# iovss 3.04218f $ **FLOATING
C73 a_6085_11542# iovss 0.41716f
C74 a_5755_7456# iovss 0.43386f
C75 a_5755_7542# iovss 3.04218f $ **FLOATING
C76 a_5425_7542# iovss 3.04218f $ **FLOATING
C77 a_5425_11542# iovss 0.41716f
C78 a_5095_7456# iovss 0.43386f
C79 a_5095_7542# iovss 3.04229f $ **FLOATING
C80 a_4765_7542# iovss 3.04218f $ **FLOATING
C81 a_4765_11542# iovss 0.41716f
C82 a_4435_7456# iovss 0.43382f
C83 a_4435_7542# iovss 3.04229f $ **FLOATING
C84 a_4105_7542# iovss 3.04218f $ **FLOATING
C85 a_4105_11542# iovss 0.41716f
C86 a_3775_7456# iovss 0.45486f
C87 a_3775_7542# iovss 3.53976f $ **FLOATING
C88 sg13g2_RCClampInverter_0.out iovss 0.24479p
C89 sg13g2_RCClampInverter_0.in iovss 0.20743p
C90 w_n124_1076# iovss 32.29903f $ **FLOATING
C91 iovdd.n0 iovss 1.37481f
C92 iovdd.n1 iovss 2.13336f
C93 iovdd.n2 iovss 0.6874f
C94 iovdd.n3 iovss 4.7379f
C95 iovdd.n4 iovss 1.37481f
C96 iovdd.n5 iovss 0.6874f
C97 iovdd.n6 iovss 1.37481f
C98 iovdd.n7 iovss 0.6874f
C99 iovdd.n8 iovss 1.37481f
C100 iovdd.n9 iovss 1.37481f
C101 iovdd.n10 iovss 1.37481f
C102 iovdd.n11 iovss 1.37481f
C103 iovdd.n12 iovss 0.6874f
C104 iovdd.n13 iovss 1.37481f
C105 iovdd.n14 iovss 0.6874f
C106 iovdd.n15 iovss 1.37481f
C107 iovdd.n16 iovss 1.37481f
C108 iovdd.n17 iovss 1.37481f
C109 iovdd.n18 iovss 1.37481f
C110 iovdd.n19 iovss 0.6874f
C111 iovdd.n20 iovss 1.37481f
C112 iovdd.n21 iovss 0.6874f
C113 iovdd.n22 iovss 1.37481f
C114 iovdd.n23 iovss 1.37481f
C115 iovdd.n24 iovss 1.37481f
C116 iovdd.n25 iovss 1.37481f
C117 iovdd.n26 iovss 0.6874f
C118 iovdd.n27 iovss 1.37481f
C119 iovdd.n28 iovss 0.6874f
C120 iovdd.n29 iovss 1.37481f
C121 iovdd.n30 iovss 1.37481f
C122 iovdd.n31 iovss 1.37481f
C123 iovdd.n32 iovss 1.37481f
C124 iovdd.n33 iovss 0.6874f
C125 iovdd.n34 iovss 1.37481f
C126 iovdd.n35 iovss 0.6874f
C127 iovdd.n36 iovss 1.37481f
C128 iovdd.n37 iovss 1.37481f
C129 iovdd.n38 iovss 1.37481f
C130 iovdd.n39 iovss 1.37481f
C131 iovdd.n40 iovss 0.6874f
C132 iovdd.n41 iovss 1.37481f
C133 iovdd.n42 iovss 0.6874f
C134 iovdd.n43 iovss 1.37481f
C135 iovdd.n44 iovss 1.37481f
C136 iovdd.n45 iovss 1.37481f
C137 iovdd.n46 iovss 1.37481f
C138 iovdd.n47 iovss 0.6874f
C139 iovdd.n48 iovss 1.37481f
C140 iovdd.n49 iovss 0.6874f
C141 iovdd.n50 iovss 1.37481f
C142 iovdd.n51 iovss 1.37481f
C143 iovdd.n52 iovss 1.37481f
C144 iovdd.n53 iovss 1.37481f
C145 iovdd.n54 iovss 0.6874f
C146 iovdd.n55 iovss 1.37481f
C147 iovdd.n56 iovss 0.6874f
C148 iovdd.n57 iovss 1.37481f
C149 iovdd.n58 iovss 1.37481f
C150 iovdd.n59 iovss 1.37481f
C151 iovdd.n60 iovss 1.37481f
C152 iovdd.n61 iovss 0.6874f
C153 iovdd.n62 iovss 1.37481f
C154 iovdd.n63 iovss 0.6874f
C155 iovdd.n64 iovss 1.37481f
C156 iovdd.n65 iovss 1.37481f
C157 iovdd.n66 iovss 1.37481f
C158 iovdd.n67 iovss 1.37481f
C159 iovdd.n68 iovss 0.6874f
C160 iovdd.n69 iovss 1.37481f
C161 iovdd.n70 iovss 0.6874f
C162 iovdd.n71 iovss 1.37481f
C163 iovdd.n72 iovss 1.37481f
C164 iovdd.n73 iovss 1.37481f
C165 iovdd.n74 iovss 1.37481f
C166 iovdd.n75 iovss 0.6874f
C167 iovdd.n76 iovss 1.37481f
C168 iovdd.n77 iovss 0.6874f
C169 iovdd.n78 iovss 1.37481f
C170 iovdd.n79 iovss 1.37481f
C171 iovdd.n80 iovss 1.37481f
C172 iovdd.n81 iovss 1.37481f
C173 iovdd.n82 iovss 0.6874f
C174 iovdd.n83 iovss 0.50474f
C175 iovdd.n84 iovss 1.56962f
C176 iovdd.n85 iovss 2.40868f
C177 iovdd.n86 iovss 4.7379f
C178 iovdd.n87 iovss 2.13336f
C179 iovdd.n88 iovss 1.37481f
C180 iovdd.n89 iovss 0.6874f
C181 iovdd.n90 iovss 0.6874f
C182 iovdd.n91 iovss 1.37481f
C183 iovdd.n92 iovss 1.37481f
C184 iovdd.n93 iovss 0.6874f
C185 iovdd.n94 iovss 0.6874f
C186 iovdd.n95 iovss 1.37481f
C187 iovdd.n96 iovss 1.37481f
C188 iovdd.n97 iovss 0.6874f
C189 iovdd.n98 iovss 0.6874f
C190 iovdd.n99 iovss 1.37481f
C191 iovdd.n100 iovss 1.37481f
C192 iovdd.n101 iovss 0.6874f
C193 iovdd.n102 iovss 0.6874f
C194 iovdd.n103 iovss 1.37481f
C195 iovdd.n104 iovss 1.37481f
C196 iovdd.n105 iovss 0.6874f
C197 iovdd.n106 iovss 0.6874f
C198 iovdd.n107 iovss 1.37481f
C199 iovdd.n108 iovss 1.37481f
C200 iovdd.n109 iovss 0.6874f
C201 iovdd.n110 iovss 0.6874f
C202 iovdd.n111 iovss 1.37481f
C203 iovdd.n112 iovss 1.37481f
C204 iovdd.n113 iovss 0.6874f
C205 iovdd.n114 iovss 0.6874f
C206 iovdd.n115 iovss 1.37481f
C207 iovdd.n116 iovss 1.37481f
C208 iovdd.n117 iovss 0.6874f
C209 iovdd.n118 iovss 0.6874f
C210 iovdd.n119 iovss 1.37481f
C211 iovdd.n120 iovss 1.37481f
C212 iovdd.n121 iovss 0.6874f
C213 iovdd.n122 iovss 0.6874f
C214 iovdd.n123 iovss 1.37481f
C215 iovdd.n124 iovss 1.37481f
C216 iovdd.n125 iovss 0.6874f
C217 iovdd.n126 iovss 0.6874f
C218 iovdd.n127 iovss 1.37481f
C219 iovdd.n128 iovss 1.37481f
C220 iovdd.n129 iovss 0.6874f
C221 iovdd.n130 iovss 0.6874f
C222 iovdd.n131 iovss 1.37481f
C223 iovdd.n132 iovss 1.37481f
C224 iovdd.n133 iovss 0.6874f
C225 iovdd.n134 iovss 0.6874f
C226 iovdd.n135 iovss 1.37481f
C227 iovdd.n136 iovss 1.37481f
C228 iovdd.n137 iovss 0.6874f
C229 iovdd.n138 iovss 0.6874f
C230 iovdd.n139 iovss 1.37481f
C231 iovdd.n140 iovss 1.37481f
C232 iovdd.n141 iovss 0.6874f
C233 iovdd.n142 iovss 0.6874f
C234 iovdd.n143 iovss 1.37481f
C235 iovdd.n144 iovss 1.37481f
C236 iovdd.n145 iovss 0.6874f
C237 iovdd.n146 iovss 0.6874f
C238 iovdd.n147 iovss 1.37481f
C239 iovdd.n148 iovss 1.37481f
C240 iovdd.n149 iovss 0.6874f
C241 iovdd.n150 iovss 0.6874f
C242 iovdd.n151 iovss 1.37481f
C243 iovdd.n152 iovss 1.37481f
C244 iovdd.n153 iovss 0.6874f
C245 iovdd.n154 iovss 0.6874f
C246 iovdd.n155 iovss 1.37481f
C247 iovdd.n156 iovss 1.37481f
C248 iovdd.n157 iovss 0.6874f
C249 iovdd.n158 iovss 0.6874f
C250 iovdd.n159 iovss 1.37481f
C251 iovdd.n160 iovss 1.37481f
C252 iovdd.n161 iovss 0.6874f
C253 iovdd.n162 iovss 0.6874f
C254 iovdd.n163 iovss 1.37481f
C255 iovdd.n164 iovss 1.37481f
C256 iovdd.n165 iovss 0.6874f
C257 iovdd.n166 iovss 0.6874f
C258 iovdd.n167 iovss 1.37481f
C259 iovdd.n168 iovss 1.37481f
C260 iovdd.n169 iovss 0.6874f
C261 iovdd.n170 iovss 0.6874f
C262 iovdd.n171 iovss 1.37481f
C263 iovdd.n172 iovss 1.37481f
C264 iovdd.n173 iovss 0.6874f
C265 iovdd.n174 iovss 0.6874f
C266 iovdd.n175 iovss 1.37481f
C267 iovdd.n176 iovss 1.37481f
C268 iovdd.n177 iovss 0.6874f
C269 iovdd.n178 iovss 0.6874f
C270 iovdd.n179 iovss 1.37481f
C271 iovdd.n180 iovss 1.37481f
C272 iovdd.n181 iovss 0.6874f
C273 iovdd.n182 iovss 0.6874f
C274 iovdd.n183 iovss 1.37481f
C275 iovdd.n184 iovss 1.37481f
C276 iovdd.n185 iovss 0.6874f
C277 iovdd.n186 iovss 2.40868f
C278 iovdd.n187 iovss 3.36336f
C279 sg13g2_RCClampInverter_0.in.t2 iovss 70.6081f
C280 sg13g2_RCClampInverter_0.in.t1 iovss 11.3294f
C281 sg13g2_RCClampInverter_0.in.n0 iovss 26.3385f
C282 sg13g2_RCClampInverter_0.in.n1 iovss 0.27382f
C283 vdd.n0 iovss 0.40047f
C284 vdd.n10 iovss 0.10622f
C285 vdd.n26 iovss 0.12017f
C286 vdd.n38 iovss 0.12017f
C287 vdd.n58 iovss 0.12017f
C288 vdd.n65 iovss 0.12017f
C289 vdd.n78 iovss 0.12017f
C290 vdd.n92 iovss 0.44943f
C291 vdd.n93 iovss 0.44943f
C292 vdd.n94 iovss 0.44943f
C293 vdd.n95 iovss 0.44943f
C294 vdd.n97 iovss 0.44943f
C295 vdd.n99 iovss 0.57209f
C296 vdd.n100 iovss 0.45767f
C297 vdd.n101 iovss 0.22472f
C298 vdd.n103 iovss 0.56722f
C299 vdd.n105 iovss 0.44943f
C300 vdd.n106 iovss 1.94272f
C301 vdd.n109 iovss 0.22472f
C302 vdd.n110 iovss 0.22472f
C303 vdd.n111 iovss 0.3945f
C304 vdd.n112 iovss 0.22472f
C305 vdd.n113 iovss 0.66802f
C306 vdd.n114 iovss 0.22472f
C307 vdd.n115 iovss 2.42995f
C308 vdd.n116 iovss 0.3945f
C309 vdd.n117 iovss 0.22472f
C310 vdd.n118 iovss 0.22472f
C311 vdd.n119 iovss 0.22472f
C312 vdd.n120 iovss 0.22472f
C313 vdd.n121 iovss 0.22472f
C314 vdd.n122 iovss 0.3945f
C315 vdd.n123 iovss 0.22472f
C316 vdd.n124 iovss 0.22472f
C317 vdd.n125 iovss 0.3945f
C318 vdd.n126 iovss 0.3945f
C319 vdd.n127 iovss 0.3945f
C320 vdd.n128 iovss 0.22472f
C321 vdd.n129 iovss 0.44943f
C322 vdd.n130 iovss 0.35861f
C323 vdd.n136 iovss 0.44943f
C324 vdd.n139 iovss 0.44943f
C325 vdd.n140 iovss 0.44943f
C326 vdd.n141 iovss 0.44943f
C327 vdd.n142 iovss 0.44943f
C328 vdd.n143 iovss 0.44943f
C329 vdd.n145 iovss 0.22472f
C330 vdd.n146 iovss 0.44943f
C331 vdd.n150 iovss 0.45767f
C332 vdd.n151 iovss 0.45767f
C333 vdd.n153 iovss 0.44943f
C334 vdd.n154 iovss 0.57209f
C335 vdd.n156 iovss 0.45767f
C336 vdd.n157 iovss 0.22472f
C337 vdd.n158 iovss 0.22472f
C338 vdd.n159 iovss 4.07113f
C339 vdd.n160 iovss 0.22472f
C340 vdd.n161 iovss 0.3945f
C341 vdd.n162 iovss 0.22472f
C342 vdd.n163 iovss 0.3945f
C343 vdd.n164 iovss 0.22472f
C344 vdd.n165 iovss 0.22472f
C345 vdd.n166 iovss 0.22472f
C346 vdd.n167 iovss 0.22472f
C347 vdd.n168 iovss 0.3945f
C348 vdd.n169 iovss 0.3945f
C349 vdd.n170 iovss 0.22472f
C350 vdd.n171 iovss 0.22472f
C351 vdd.n172 iovss 0.22472f
C352 vdd.n173 iovss 0.22472f
C353 vdd.n174 iovss 0.22472f
C354 vdd.n175 iovss 0.3945f
C355 vdd.n176 iovss 0.29588f
C356 vdd.n177 iovss 0.22472f
C357 vdd.n178 iovss 0.22472f
C358 vdd.n180 iovss 0.44943f
C359 vdd.n181 iovss 0.22472f
C360 vdd.n182 iovss 0.22472f
C361 vdd.n183 iovss 0.37827f
C362 vdd.n184 iovss 0.50437f
C363 vdd.n185 iovss 0.50437f
C364 vdd.n186 iovss 0.22472f
C365 vdd.n187 iovss 0.44943f
C366 vdd.n190 iovss 0.44943f
C367 vdd.n191 iovss 0.44943f
C368 vdd.n192 iovss 0.44943f
C369 vdd.n193 iovss 0.44943f
C370 vdd.n194 iovss 0.44943f
C371 vdd.n196 iovss 0.44943f
C372 vdd.n197 iovss 0.57209f
C373 vdd.n198 iovss 0.45767f
C374 vdd.n201 iovss 0.45767f
C375 vdd.n202 iovss 0.22472f
C376 vdd.n203 iovss 0.44943f
C377 vdd.n207 iovss 0.45767f
C378 vdd.n210 iovss 0.22472f
C379 vdd.n211 iovss 0.22472f
C380 vdd.n212 iovss 0.11318f
C381 vdd.t0 iovss 7.475f
C382 vdd.n266 iovss 0.49034f
C383 vdd.n268 iovss 15.3572f
C384 vdd.n269 iovss 34.1576f
C385 vdd.n270 iovss 0.57733f
C386 vdd.n271 iovss 0.22472f
C387 vdd.n272 iovss 0.50437f
C388 vdd.n273 iovss 0.22472f
C389 vdd.n274 iovss 0.22472f
C390 vdd.n275 iovss 0.50437f
C391 vdd.n276 iovss 0.50437f
C392 vdd.n277 iovss 0.22472f
C393 vdd.n278 iovss 0.22472f
C394 vdd.n279 iovss 0.22472f
C395 vdd.n280 iovss 0.22472f
C396 vdd.n281 iovss 0.22472f
C397 vdd.n282 iovss 0.22472f
C398 vdd.n283 iovss 0.50437f
C399 vdd.n284 iovss 0.50437f
C400 vdd.n285 iovss 0.50437f
C401 vdd.n286 iovss 0.22472f
C402 vdd.n287 iovss 0.50437f
C403 vdd.n288 iovss 0.40012f
C404 vdd.n289 iovss 0.37827f
C405 vdd.n290 iovss 0.33708f
C406 vdd.n291 iovss 0.2304f
C407 vdd.n292 iovss 1.34262f
C408 vdd.n293 iovss 0.22472f
C409 vdd.n294 iovss 0.22472f
C410 vdd.n295 iovss 0.22472f
C411 vdd.n296 iovss 0.22472f
C412 vdd.n297 iovss 0.50437f
C413 vdd.n298 iovss 0.50437f
C414 vdd.n299 iovss 0.22472f
C415 vdd.n300 iovss 0.22472f
C416 vdd.n301 iovss 0.22472f
C417 vdd.n302 iovss 0.50437f
C418 vdd.n303 iovss 0.50437f
C419 vdd.n304 iovss 0.22472f
C420 vdd.n305 iovss 0.22472f
C421 vdd.n307 iovss 0.44943f
C422 vdd.n309 iovss 0.45767f
C423 vdd.n310 iovss 0.44943f
C424 vdd.n311 iovss 2.2835f
C425 vdd.n312 iovss 0.29681f
C426 vdd.n313 iovss 0.44943f
C427 vdd.n314 iovss 0.22472f
C428 vdd.n315 iovss 0.22472f
C429 vdd.n316 iovss 0.22472f
C430 vdd.n317 iovss 0.22472f
C431 vdd.n318 iovss 0.50437f
C432 vdd.n319 iovss 0.22472f
C433 vdd.n320 iovss 0.50437f
C434 vdd.n321 iovss 0.50437f
C435 vdd.n322 iovss 0.22472f
C436 vdd.n323 iovss 0.22472f
C437 vdd.n324 iovss 0.44943f
C438 vdd.n325 iovss 0.40047f
C439 vdd.n326 iovss 0.44943f
C440 vdd.n327 iovss 0.45767f
C441 vdd.n329 iovss 4.70203f
C442 vdd.n330 iovss 0.35955f
C443 vdd.n331 iovss 0.29681f
C444 vdd.n332 iovss 0.44943f
C445 vdd.n333 iovss 0.22472f
C446 vdd.n334 iovss 0.22472f
C447 vdd.n335 iovss 0.3945f
C448 vdd.n336 iovss 0.3945f
C449 vdd.n337 iovss 0.22472f
C450 vdd.n338 iovss 0.22472f
C451 vdd.n339 iovss 0.44943f
C452 vdd.n343 iovss 0.45767f
C453 vdd.n345 iovss 0.45767f
C454 vdd.n347 iovss 2.35501f
C455 vdd.n349 iovss 0.45767f
C456 vdd.n350 iovss 0.44943f
C457 vdd.n351 iovss 0.40047f
C458 vdd.n369 iovss 0.12017f
C459 vdd.n376 iovss 0.12017f
C460 vdd.n381 iovss 0.12017f
C461 vdd.n388 iovss 0.12017f
C462 vdd.n397 iovss 0.12017f
C463 vdd.n404 iovss 0.12017f
C464 vdd.n407 iovss 0.11214f
C465 vdd.n433 iovss 0.12017f
C466 vdd.n487 iovss 0.12017f
C467 vdd.n494 iovss 0.12017f
C468 vdd.n500 iovss 0.12017f
C469 vdd.n556 iovss 17.5508f
C470 vdd.n584 iovss 0.12017f
C471 vdd.n591 iovss 0.12017f
C472 vdd.n643 iovss 0.12017f
C473 vdd.n662 iovss 17.0485f
C474 vdd.n686 iovss 0.12017f
C475 vdd.n724 iovss 0.12017f
C476 vdd.n736 iovss 0.12017f
C477 vdd.n763 iovss 0.12017f
C478 vdd.n778 iovss 0.17924f
C479 vdd.n784 iovss 16.6116f
C480 sg13g2_RCClampInverter_0.out.t66 iovss 0.9055f
C481 sg13g2_RCClampInverter_0.out.t109 iovss 0.51153f
C482 sg13g2_RCClampInverter_0.out.n0 iovss 0.11866f
C483 sg13g2_RCClampInverter_0.out.t70 iovss 0.9055f
C484 sg13g2_RCClampInverter_0.out.t85 iovss 0.51153f
C485 sg13g2_RCClampInverter_0.out.n2 iovss 0.36603f
C486 sg13g2_RCClampInverter_0.out.t88 iovss 0.9055f
C487 sg13g2_RCClampInverter_0.out.t32 iovss 0.51153f
C488 sg13g2_RCClampInverter_0.out.n4 iovss 0.2025f
C489 sg13g2_RCClampInverter_0.out.t37 iovss 0.9055f
C490 sg13g2_RCClampInverter_0.out.t99 iovss 0.51153f
C491 sg13g2_RCClampInverter_0.out.n6 iovss 0.2025f
C492 sg13g2_RCClampInverter_0.out.t51 iovss 0.9055f
C493 sg13g2_RCClampInverter_0.out.t68 iovss 0.51153f
C494 sg13g2_RCClampInverter_0.out.n8 iovss 0.2025f
C495 sg13g2_RCClampInverter_0.out.t60 iovss 0.9055f
C496 sg13g2_RCClampInverter_0.out.t103 iovss 0.51153f
C497 sg13g2_RCClampInverter_0.out.n10 iovss 0.2025f
C498 sg13g2_RCClampInverter_0.out.t75 iovss 0.9055f
C499 sg13g2_RCClampInverter_0.out.t89 iovss 0.51153f
C500 sg13g2_RCClampInverter_0.out.n12 iovss 0.2025f
C501 sg13g2_RCClampInverter_0.out.t98 iovss 0.9055f
C502 sg13g2_RCClampInverter_0.out.t47 iovss 0.51153f
C503 sg13g2_RCClampInverter_0.out.n14 iovss 0.2025f
C504 sg13g2_RCClampInverter_0.out.t58 iovss 0.9055f
C505 sg13g2_RCClampInverter_0.out.t72 iovss 0.51153f
C506 sg13g2_RCClampInverter_0.out.n16 iovss 0.2025f
C507 sg13g2_RCClampInverter_0.out.t53 iovss 0.9055f
C508 sg13g2_RCClampInverter_0.out.t69 iovss 0.51153f
C509 sg13g2_RCClampInverter_0.out.n18 iovss 0.2025f
C510 sg13g2_RCClampInverter_0.out.t45 iovss 0.9055f
C511 sg13g2_RCClampInverter_0.out.t106 iovss 0.51153f
C512 sg13g2_RCClampInverter_0.out.n20 iovss 0.2025f
C513 sg13g2_RCClampInverter_0.out.t36 iovss 0.9055f
C514 sg13g2_RCClampInverter_0.out.t50 iovss 0.51153f
C515 sg13g2_RCClampInverter_0.out.n22 iovss 0.2025f
C516 sg13g2_RCClampInverter_0.out.t67 iovss 0.9055f
C517 sg13g2_RCClampInverter_0.out.t110 iovss 0.51153f
C518 sg13g2_RCClampInverter_0.out.n24 iovss 0.2025f
C519 sg13g2_RCClampInverter_0.out.t56 iovss 0.9055f
C520 sg13g2_RCClampInverter_0.out.t102 iovss 0.51153f
C521 sg13g2_RCClampInverter_0.out.n26 iovss 0.2025f
C522 sg13g2_RCClampInverter_0.out.t33 iovss 0.9055f
C523 sg13g2_RCClampInverter_0.out.t49 iovss 0.51153f
C524 sg13g2_RCClampInverter_0.out.n28 iovss 0.2025f
C525 sg13g2_RCClampInverter_0.out.t34 iovss 0.9055f
C526 sg13g2_RCClampInverter_0.out.t105 iovss 0.51153f
C527 sg13g2_RCClampInverter_0.out.n30 iovss 0.2025f
C528 sg13g2_RCClampInverter_0.out.t86 iovss 0.9055f
C529 sg13g2_RCClampInverter_0.out.t96 iovss 0.51153f
C530 sg13g2_RCClampInverter_0.out.n32 iovss 0.2025f
C531 sg13g2_RCClampInverter_0.out.t41 iovss 0.9055f
C532 sg13g2_RCClampInverter_0.out.t55 iovss 0.51153f
C533 sg13g2_RCClampInverter_0.out.n34 iovss 0.2025f
C534 sg13g2_RCClampInverter_0.out.t65 iovss 0.9055f
C535 sg13g2_RCClampInverter_0.out.t82 iovss 0.51153f
C536 sg13g2_RCClampInverter_0.out.n36 iovss 0.2025f
C537 sg13g2_RCClampInverter_0.out.t62 iovss 0.9055f
C538 sg13g2_RCClampInverter_0.out.t78 iovss 0.51153f
C539 sg13g2_RCClampInverter_0.out.n38 iovss 0.2025f
C540 sg13g2_RCClampInverter_0.out.t54 iovss 0.9055f
C541 sg13g2_RCClampInverter_0.out.t108 iovss 0.51153f
C542 sg13g2_RCClampInverter_0.out.n40 iovss 0.2025f
C543 sg13g2_RCClampInverter_0.out.t46 iovss 0.9055f
C544 sg13g2_RCClampInverter_0.out.t61 iovss 0.51153f
C545 sg13g2_RCClampInverter_0.out.n42 iovss 0.2025f
C546 sg13g2_RCClampInverter_0.out.t77 iovss 0.9055f
C547 sg13g2_RCClampInverter_0.out.t115 iovss 0.51153f
C548 sg13g2_RCClampInverter_0.out.n44 iovss 0.2025f
C549 sg13g2_RCClampInverter_0.out.t31 iovss 0.9055f
C550 sg13g2_RCClampInverter_0.out.t104 iovss 0.51153f
C551 sg13g2_RCClampInverter_0.out.n46 iovss 0.2025f
C552 sg13g2_RCClampInverter_0.out.t42 iovss 0.9055f
C553 sg13g2_RCClampInverter_0.out.t57 iovss 0.51153f
C554 sg13g2_RCClampInverter_0.out.n48 iovss 0.2025f
C555 sg13g2_RCClampInverter_0.out.t48 iovss 0.9055f
C556 sg13g2_RCClampInverter_0.out.t101 iovss 0.51153f
C557 sg13g2_RCClampInverter_0.out.n50 iovss 0.2025f
C558 sg13g2_RCClampInverter_0.out.t63 iovss 0.9055f
C559 sg13g2_RCClampInverter_0.out.t80 iovss 0.51153f
C560 sg13g2_RCClampInverter_0.out.n52 iovss 0.2025f
C561 sg13g2_RCClampInverter_0.out.t90 iovss 0.9055f
C562 sg13g2_RCClampInverter_0.out.t35 iovss 0.51153f
C563 sg13g2_RCClampInverter_0.out.n54 iovss 0.2025f
C564 sg13g2_RCClampInverter_0.out.t87 iovss 0.9055f
C565 sg13g2_RCClampInverter_0.out.t97 iovss 0.51153f
C566 sg13g2_RCClampInverter_0.out.n56 iovss 0.2025f
C567 sg13g2_RCClampInverter_0.out.t43 iovss 0.9055f
C568 sg13g2_RCClampInverter_0.out.t59 iovss 0.51153f
C569 sg13g2_RCClampInverter_0.out.n58 iovss 0.2025f
C570 sg13g2_RCClampInverter_0.out.t74 iovss 0.9055f
C571 sg13g2_RCClampInverter_0.out.t112 iovss 0.51153f
C572 sg13g2_RCClampInverter_0.out.n60 iovss 0.2025f
C573 sg13g2_RCClampInverter_0.out.t92 iovss 0.9055f
C574 sg13g2_RCClampInverter_0.out.t39 iovss 0.51153f
C575 sg13g2_RCClampInverter_0.out.n62 iovss 0.2025f
C576 sg13g2_RCClampInverter_0.out.t93 iovss 0.9055f
C577 sg13g2_RCClampInverter_0.out.t40 iovss 0.51153f
C578 sg13g2_RCClampInverter_0.out.n64 iovss 0.2025f
C579 sg13g2_RCClampInverter_0.out.t44 iovss 0.9055f
C580 sg13g2_RCClampInverter_0.out.t100 iovss 0.51153f
C581 sg13g2_RCClampInverter_0.out.n66 iovss 0.2025f
C582 sg13g2_RCClampInverter_0.out.t79 iovss 0.9055f
C583 sg13g2_RCClampInverter_0.out.t116 iovss 0.51153f
C584 sg13g2_RCClampInverter_0.out.n68 iovss 0.2025f
C585 sg13g2_RCClampInverter_0.out.t83 iovss 0.9055f
C586 sg13g2_RCClampInverter_0.out.t94 iovss 0.51153f
C587 sg13g2_RCClampInverter_0.out.n70 iovss 0.2025f
C588 sg13g2_RCClampInverter_0.out.t84 iovss 0.9055f
C589 sg13g2_RCClampInverter_0.out.t95 iovss 0.51153f
C590 sg13g2_RCClampInverter_0.out.n72 iovss 0.2025f
C591 sg13g2_RCClampInverter_0.out.t71 iovss 0.9055f
C592 sg13g2_RCClampInverter_0.out.t111 iovss 0.51153f
C593 sg13g2_RCClampInverter_0.out.n74 iovss 0.2025f
C594 sg13g2_RCClampInverter_0.out.t64 iovss 0.9055f
C595 sg13g2_RCClampInverter_0.out.t81 iovss 0.51153f
C596 sg13g2_RCClampInverter_0.out.n76 iovss 0.2025f
C597 sg13g2_RCClampInverter_0.out.t91 iovss 0.9055f
C598 sg13g2_RCClampInverter_0.out.t38 iovss 0.51153f
C599 sg13g2_RCClampInverter_0.out.n78 iovss 0.2025f
C600 sg13g2_RCClampInverter_0.out.t52 iovss 0.9055f
C601 sg13g2_RCClampInverter_0.out.t107 iovss 0.51153f
C602 sg13g2_RCClampInverter_0.out.n80 iovss 0.2025f
C603 sg13g2_RCClampInverter_0.out.t73 iovss 0.9055f
C604 sg13g2_RCClampInverter_0.out.t113 iovss 0.51153f
C605 sg13g2_RCClampInverter_0.out.n82 iovss 0.2025f
C606 sg13g2_RCClampInverter_0.out.t76 iovss 0.9055f
C607 sg13g2_RCClampInverter_0.out.t114 iovss 0.51153f
C608 sg13g2_RCClampInverter_0.out.n84 iovss 0.22436f
C609 sg13g2_RCClampInverter_0.out.t17 iovss 0.3917f
C610 sg13g2_RCClampInverter_0.out.t19 iovss 0.38065f
C611 sg13g2_RCClampInverter_0.out.n86 iovss 2.25104f
C612 sg13g2_RCClampInverter_0.out.t20 iovss 0.38065f
C613 sg13g2_RCClampInverter_0.out.n87 iovss 1.42996f
C614 sg13g2_RCClampInverter_0.out.t24 iovss 0.38065f
C615 sg13g2_RCClampInverter_0.out.n88 iovss 1.42996f
C616 sg13g2_RCClampInverter_0.out.t28 iovss 0.38065f
C617 sg13g2_RCClampInverter_0.out.n89 iovss 1.42996f
C618 sg13g2_RCClampInverter_0.out.t29 iovss 0.38065f
C619 sg13g2_RCClampInverter_0.out.n90 iovss 1.42996f
C620 sg13g2_RCClampInverter_0.out.t14 iovss 0.38065f
C621 sg13g2_RCClampInverter_0.out.n91 iovss 1.42996f
C622 sg13g2_RCClampInverter_0.out.t13 iovss 0.38065f
C623 sg13g2_RCClampInverter_0.out.n92 iovss 1.42996f
C624 sg13g2_RCClampInverter_0.out.t23 iovss 0.38065f
C625 sg13g2_RCClampInverter_0.out.n93 iovss 1.42996f
C626 sg13g2_RCClampInverter_0.out.t22 iovss 0.38065f
C627 sg13g2_RCClampInverter_0.out.n94 iovss 1.42996f
C628 sg13g2_RCClampInverter_0.out.t11 iovss 0.38065f
C629 sg13g2_RCClampInverter_0.out.n95 iovss 1.42996f
C630 sg13g2_RCClampInverter_0.out.t10 iovss 0.38065f
C631 sg13g2_RCClampInverter_0.out.n96 iovss 1.42996f
C632 sg13g2_RCClampInverter_0.out.t12 iovss 0.38065f
C633 sg13g2_RCClampInverter_0.out.n97 iovss 1.42996f
C634 sg13g2_RCClampInverter_0.out.t18 iovss 0.38065f
C635 sg13g2_RCClampInverter_0.out.n98 iovss 1.42996f
C636 sg13g2_RCClampInverter_0.out.t9 iovss 0.38065f
C637 sg13g2_RCClampInverter_0.out.n99 iovss 1.42996f
C638 sg13g2_RCClampInverter_0.out.t8 iovss 0.38065f
C639 sg13g2_RCClampInverter_0.out.n100 iovss 1.42996f
C640 sg13g2_RCClampInverter_0.out.t7 iovss 0.38065f
C641 sg13g2_RCClampInverter_0.out.n101 iovss 1.42996f
C642 sg13g2_RCClampInverter_0.out.t26 iovss 0.38065f
C643 sg13g2_RCClampInverter_0.out.n102 iovss 1.42996f
C644 sg13g2_RCClampInverter_0.out.t25 iovss 0.38065f
C645 sg13g2_RCClampInverter_0.out.n103 iovss 1.42996f
C646 sg13g2_RCClampInverter_0.out.t30 iovss 0.38065f
C647 sg13g2_RCClampInverter_0.out.n104 iovss 1.42996f
C648 sg13g2_RCClampInverter_0.out.t27 iovss 0.38065f
C649 sg13g2_RCClampInverter_0.out.n105 iovss 1.42996f
C650 sg13g2_RCClampInverter_0.out.t21 iovss 0.38065f
C651 sg13g2_RCClampInverter_0.out.n106 iovss 1.42996f
C652 sg13g2_RCClampInverter_0.out.t16 iovss 0.38065f
C653 sg13g2_RCClampInverter_0.out.n107 iovss 1.42996f
C654 sg13g2_RCClampInverter_0.out.t15 iovss 0.38065f
C655 sg13g2_RCClampInverter_0.out.n108 iovss 1.42996f
C656 sg13g2_RCClampInverter_0.out.t6 iovss 0.38066f
C657 sg13g2_RCClampInverter_0.out.n109 iovss 12.0539f
C658 sg13g2_RCClampInverter_0.out.t4 iovss 0.5001f
C659 sg13g2_RCClampInverter_0.out.t2 iovss 0.5001f
C660 sg13g2_RCClampInverter_0.out.t0 iovss 0.5001f
C661 sg13g2_RCClampInverter_0.out.n110 iovss 15.0457f
C662 sg13g2_RCClampInverter_0.out.t1 iovss 0.5001f
C663 sg13g2_RCClampInverter_0.out.t3 iovss 0.5001f
C664 sg13g2_RCClampInverter_0.out.t5 iovss 0.49998f
C665 sg13g2_RCClampInverter_0.out.n111 iovss 5.58445f
.ends

