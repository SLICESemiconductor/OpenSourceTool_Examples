* NGSPICE file created from sg13g2_IOPadInOut30mA_flat.ext - technology: ihp-sg13g2

.subckt sg13g2_IOPadInOut30mA_flat p2c c2p_en c2p pad vdd iovdd iovss
X0 vdd a_12038_31490# p2c vdd sg13_lv_pmos ad=1.615p pd=10.18u as=1.615p ps=10.18u w=4.75u l=0.13u
X1 sg13g2_GateDecode_0.pgate iovdd dpantenna l=0.78u w=0.78u
X2 iovdd sg13g2_GateDecode_0.pgate pad iovdd sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X3 iovdd sg13g2_GateDecode_0.pgate pad iovdd sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X4 iovss sg13g2_GateDecode_0.ngate pad iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X5 pad sg13g2_GateDecode_0.pgate iovdd iovdd sg13_hv_pmos ad=3.9294p pd=7.84u as=3.1302p ps=14.26u w=6.66u l=0.6u
X6 iovdd sg13g2_GateDecode_0.pgate pad iovdd sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X7 pad sg13g2_GateDecode_0.pgate iovdd iovdd sg13_hv_pmos ad=4.9284p pd=14.8u as=2.1312p ps=7.3u w=6.66u l=0.6u
X8 iovss a_12038_31490# p2c iovss sg13_lv_nmos ad=0.935p pd=6.18u as=0.935p ps=6.18u w=2.75u l=0.13u
X9 iovdd sg13g2_GateDecode_0.pgate pad iovdd sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X10 iovss pad dantenna l=1.26u w=27.78u
X11 pad sg13g2_GateDecode_0.ngate iovss iovss sg13_hv_nmos ad=3.256p pd=10.28u as=1.408p ps=5.04u w=4.4u l=0.6u
X12 pad sg13g2_GateDecode_0.ngate iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X13 iovss sg13g2_GateDecode_0.ngate pad iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X14 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq c2p_en a_4230_33842# iovss sg13_lv_nmos ad=1.4148p pd=8.58u as=0.7467p ps=4.31u w=3.93u l=0.13u
X15 iovss sg13g2_LevelDown_0.sg13g2_SecondaryProtection_0.core dantenna l=3.1u w=0.64u
X16 pad sg13g2_GateDecode_0.pgate iovdd iovdd sg13_hv_pmos ad=3.9294p pd=7.84u as=3.1302p ps=14.26u w=6.66u l=0.6u
X17 iovdd sg13g2_GateDecode_0.pgate pad iovdd sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X18 iovdd sg13g2_GateDecode_0.pgate pad iovdd sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X19 iovss sg13g2_GateDecode_0.ngate pad iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X20 pad sg13g2_GateDecode_0.pgate iovdd iovdd sg13_hv_pmos ad=4.9284p pd=14.8u as=2.1312p ps=7.3u w=6.66u l=0.6u
X21 iovdd sg13g2_GateDecode_0.pgate pad iovdd sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X22 iovss sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq iovss sg13_lv_nmos ad=1.4148p pd=8.58u as=0.7467p ps=4.31u w=3.93u l=0.13u
X23 a_12038_31490# sg13g2_LevelDown_0.sg13g2_SecondaryProtection_0.core vdd vdd sg13_hv_pmos ad=1.581p pd=9.98u as=1.581p ps=9.98u w=4.65u l=0.45u
X24 a_3724_30170# sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq iovss iovss sg13_hv_nmos ad=0.646p pd=4.48u as=0.361p ps=2.28u w=1.9u l=0.45u
X25 iovdd a_3724_30170# a_3656_30206# iovdd sg13_hv_pmos ad=57f pd=0.68u as=0.102p ps=1.28u w=0.3u l=0.45u
X26 sg13g2_GateDecode_0.ngate a_3724_30170# iovdd iovdd sg13_hv_pmos ad=1.326p pd=8.48u as=1.326p ps=8.48u w=3.9u l=0.45u
X27 iovdd sg13g2_GateDecode_0.pgate pad iovdd sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X28 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq c2p vdd vdd sg13_lv_pmos ad=0.8379p pd=4.79u as=1.4994p ps=9.5u w=4.41u l=0.13u
X29 pad sg13g2_GateDecode_0.pgate iovdd iovdd sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X30 pad sg13g2_GateDecode_0.ngate iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X31 iovss sg13g2_GateDecode_0.ngate pad iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X32 pad sg13g2_GateDecode_0.ngate iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X33 a_4426_30170# a_4358_30206# iovdd iovdd sg13_hv_pmos ad=0.102p pd=1.28u as=57f ps=0.68u w=0.3u l=0.45u
X34 iovdd sg13g2_GateDecode_0.pgate pad iovdd sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X35 a_3750_34876# c2p vdd vdd sg13_lv_pmos ad=0.8379p pd=4.79u as=1.4994p ps=9.5u w=4.41u l=0.13u
X36 pad sg13g2_GateDecode_0.pgate iovdd iovdd sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X37 pad sg13g2_GateDecode_0.pgate iovdd iovdd sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X38 pad sg13g2_GateDecode_0.ngate iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=2.068p ps=9.74u w=4.4u l=0.6u
X39 pad sg13g2_GateDecode_0.ngate iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X40 sg13g2_GateDecode_0.ngate a_3724_30170# iovss iovss sg13_hv_nmos ad=0.646p pd=4.48u as=0.646p ps=4.48u w=1.9u l=0.45u
X41 pad sg13g2_GateDecode_0.pgate iovdd iovdd sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X42 iovdd sg13g2_GateDecode_0.pgate pad iovdd sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X43 vdd sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq a_4358_31526# vdd sg13_lv_pmos ad=1.615p pd=10.18u as=1.615p ps=10.18u w=4.75u l=0.13u
X44 iovss sg13g2_GateDecode_0.ngate dantenna l=0.78u w=0.78u
X45 iovss a_4358_31526# a_4358_30206# iovss sg13_hv_nmos ad=0.361p pd=2.28u as=0.646p ps=4.48u w=1.9u l=0.45u
X46 pad iovdd dpantenna l=1.26u w=27.78u
X47 sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq c2p_en iovss iovss sg13_lv_nmos ad=1.3362p pd=8.54u as=1.3362p ps=8.54u w=3.93u l=0.13u
X48 iovss sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq a_4358_31526# iovss sg13_lv_nmos ad=0.935p pd=6.18u as=0.935p ps=6.18u w=2.75u l=0.13u
X49 pad sg13g2_GateDecode_0.pgate iovdd iovdd sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X50 pad sg13g2_GateDecode_0.pgate iovdd iovdd sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X51 iovss sg13g2_GateDecode_0.ngate pad iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X52 iovdd sg13g2_GateDecode_0.pgate pad iovdd sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X53 pad sg13g2_GateDecode_0.pgate iovdd iovdd sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X54 vdd c2p_en sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq vdd sg13_lv_pmos ad=1.5876p pd=9.54u as=0.8379p ps=4.79u w=4.41u l=0.13u
X55 sg13g2_LevelDown_0.sg13g2_SecondaryProtection_0.core pad iovss rppd l=2u w=1u
X56 iovss sg13g2_GateDecode_0.ngate pad iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X57 sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq a_3750_34876# vdd sg13_lv_pmos ad=1.5876p pd=9.54u as=0.8379p ps=4.79u w=4.41u l=0.13u
X58 a_3724_30170# a_3656_30206# iovdd iovdd sg13_hv_pmos ad=0.102p pd=1.28u as=57f ps=0.68u w=0.3u l=0.45u
X59 iovss sg13g2_GateDecode_0.ngate pad iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X60 pad sg13g2_GateDecode_0.pgate iovdd iovdd sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X61 pad sg13g2_GateDecode_0.pgate iovdd iovdd sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X62 pad iovdd dpantenna l=1.26u w=27.78u
X63 iovdd sg13g2_GateDecode_0.pgate pad iovdd sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X64 sg13g2_GateDecode_0.pgate a_4426_30170# iovdd iovdd sg13_hv_pmos ad=1.326p pd=8.48u as=1.326p ps=8.48u w=3.9u l=0.45u
X65 pad sg13g2_GateDecode_0.ngate iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X66 vdd sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq a_3656_31526# vdd sg13_lv_pmos ad=1.615p pd=10.18u as=1.615p ps=10.18u w=4.75u l=0.13u
X67 iovss pad dantenna l=1.26u w=27.78u
X68 a_4230_33842# c2p iovss iovss sg13_lv_nmos ad=0.7467p pd=4.31u as=1.3362p ps=8.54u w=3.93u l=0.13u
X69 iovss a_3656_31526# a_3656_30206# iovss sg13_hv_nmos ad=0.361p pd=2.28u as=0.646p ps=4.48u w=1.9u l=0.45u
X70 sg13g2_LevelDown_0.sg13g2_SecondaryProtection_0.core iovdd dpantenna l=0.64u w=4.98u
X71 iovdd sg13g2_GateDecode_0.pgate pad iovdd sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X72 pad sg13g2_GateDecode_0.pgate iovdd iovdd sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X73 pad sg13g2_GateDecode_0.pgate iovdd iovdd sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X74 iovdd sg13g2_GateDecode_0.pgate pad iovdd sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X75 iovss sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq a_3656_31526# iovss sg13_lv_nmos ad=0.935p pd=6.18u as=0.935p ps=6.18u w=2.75u l=0.13u
X76 a_4426_30170# sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq iovss iovss sg13_hv_nmos ad=0.646p pd=4.48u as=0.361p ps=2.28u w=1.9u l=0.45u
X77 iovdd a_4426_30170# a_4358_30206# iovdd sg13_hv_pmos ad=57f pd=0.68u as=0.102p ps=1.28u w=0.3u l=0.45u
X78 pad sg13g2_GateDecode_0.ngate iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X79 sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq c2p iovss iovss sg13_lv_nmos ad=0.7467p pd=4.31u as=1.3362p ps=8.54u w=3.93u l=0.13u
X80 pad sg13g2_GateDecode_0.pgate iovdd iovdd sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X81 sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq c2p_en vdd vdd sg13_lv_pmos ad=1.4994p pd=9.5u as=1.4994p ps=9.5u w=4.41u l=0.13u
X82 a_12038_31490# sg13g2_LevelDown_0.sg13g2_SecondaryProtection_0.core iovss iovss sg13_hv_nmos ad=0.901p pd=5.98u as=0.901p ps=5.98u w=2.65u l=0.45u
X83 sg13g2_GateDecode_0.pgate a_4426_30170# iovss iovss sg13_hv_nmos ad=0.646p pd=4.48u as=0.646p ps=4.48u w=1.9u l=0.45u
C0 p2c a_12038_31490# 0.25311f
C1 sg13g2_LevelDown_0.sg13g2_SecondaryProtection_0.core vdd 0.51442f
C2 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq a_4426_30170# 0.1286f
C3 p2c vdd 2.6001f
C4 sg13g2_LevelDown_0.sg13g2_SecondaryProtection_0.core p2c 0.10336f
C5 a_4358_31526# sg13g2_GateDecode_0.ngate 0.42695f
C6 sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq a_3724_30170# 0.1286f
C7 c2p sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq 0.56766f
C8 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq c2p 0.43902f
C9 pad sg13g2_GateDecode_0.pgate 16.798f
C10 c2p_en c2p 0.53273f
C11 sg13g2_LevelDown_0.sg13g2_SecondaryProtection_0.core iovdd 1.37355f
C12 a_4358_31526# a_4358_30206# 0.15491f
C13 sg13g2_GateDecode_0.ngate sg13g2_GateDecode_0.pgate 1.51739f
C14 c2p_en sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq 1.6012f
C15 c2p_en sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq 1.59673f
C16 a_3724_30170# sg13g2_GateDecode_0.ngate 0.142f
C17 pad sg13g2_GateDecode_0.ngate 6.46854f
C18 iovdd sg13g2_GateDecode_0.pgate 46.53503f
C19 sg13g2_DCNDiode_0.guard pad 7.46684f
C20 a_4426_30170# sg13g2_GateDecode_0.pgate 0.142f
C21 a_3724_30170# a_3656_30206# 0.37106f
C22 a_4358_31526# sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq 0.99584f
C23 sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq a_3656_31526# 0.99218f
C24 c2p sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq 0.65338f
C25 iovdd a_3724_30170# 0.84924f
C26 pad iovdd 47.63779f
C27 vdd a_3656_31526# 0.79605f
C28 c2p vdd 1.52081f
C29 sg13g2_DCNDiode_0.guard sg13g2_GateDecode_0.ngate 3.6775f
C30 sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq 1.30685f
C31 sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq vdd 1.00261f
C32 iovdd sg13g2_GateDecode_0.ngate 6.54248f
C33 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq vdd 2.11533f
C34 iovdd a_3656_30206# 0.30461f
C35 a_4426_30170# iovdd 0.84126f
C36 c2p_en vdd 1.46533f
C37 a_4358_30206# sg13g2_GateDecode_0.ngate 0.59735f
C38 a_4358_31526# sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq 0.30586f
C39 a_4358_31526# vdd 0.81747f
C40 a_3656_31526# a_3656_30206# 0.15491f
C41 a_4358_30206# iovdd 0.28407f
C42 a_4426_30170# a_4358_30206# 0.37106f
C43 a_12038_31490# vdd 1.10866f
C44 sg13g2_LevelDown_0.sg13g2_SecondaryProtection_0.core a_12038_31490# 0.31408f
C45 sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq vdd 1.87035f
C46 pad iovss 0.1328p
C47 p2c iovss 2.10209f
C48 c2p_en iovss 2.18641f
C49 c2p iovss 2.43746f
C50 iovdd iovss 0.14212p
C51 vdd iovss 0.24618p
C52 a_12137_28308# iovss 0.47362f $ **FLOATING
C53 sg13g2_GateDecode_0.pgate iovss 28.34186f
C54 a_4358_30206# iovss 0.23648f
C55 sg13g2_GateDecode_0.ngate iovss 47.00961f
C56 a_3656_30206# iovss 0.45339f
C57 a_4426_30170# iovss 1.28302f
C58 a_3724_30170# iovss 1.27692f
C59 sg13g2_LevelDown_0.sg13g2_SecondaryProtection_0.core iovss 6.27806f
C60 a_4358_31526# iovss 1.33907f
C61 a_3656_31526# iovss 1.89714f
C62 a_12038_31490# iovss 1.36953f
C63 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq iovss 3.02598f
C64 sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq iovss 2.73965f
C65 sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq iovss 1.32815f
C66 sg13g2_DCNDiode_0.guard iovss 53.69175f $ **FLOATING
.ends

