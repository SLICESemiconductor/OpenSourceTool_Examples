* NGSPICE file created from sg13g2_IOPadIOVdd_flat.ext - technology: ihp-sg13g2

.subckt sg13g2_IOPadIOVdd_flat iovdd vdd vss iovss
X0 iovss sg13g2_Clamp_N43N43D4R_0.gate.t31 iovdd.t66 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X1 iovdd.t80 sg13g2_Clamp_N43N43D4R_0.gate.t32 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X2 iovdd.t68 sg13g2_Clamp_N43N43D4R_0.gate.t33 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X3 iovdd.t131 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t9 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X4 sg13g2_Clamp_N43N43D4R_0.gate.t30 sg13g2_RCClampResistor_0.pin2.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=1.71p ps=9.38u w=9u l=0.5u
X5 iovss sg13g2_Clamp_N43N43D4R_0.gate.t34 iovdd.t38 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X6 iovss sg13g2_Clamp_N43N43D4R_0.gate.t35 iovdd.t74 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X7 iovss sg13g2_Clamp_N43N43D4R_0.gate.t36 iovdd.t37 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X8 iovdd.t115 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t21 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X9 sg13g2_Clamp_N43N43D4R_0.gate.t29 sg13g2_RCClampResistor_0.pin2.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=1.71p ps=9.38u w=9u l=0.5u
X10 iovss sg13g2_Clamp_N43N43D4R_0.gate.t37 iovdd.t35 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X11 iovss sg13g2_Clamp_N43N43D4R_0.gate.t38 iovdd.t33 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X12 iovss sg13g2_Clamp_N43N43D4R_0.gate.t39 iovdd.t87 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X13 iovdd.t87 sg13g2_Clamp_N43N43D4R_0.gate.t40 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X14 iovss sg13g2_Clamp_N43N43D4R_0.gate.t41 iovdd.t86 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X15 iovdd.t62 sg13g2_Clamp_N43N43D4R_0.gate.t42 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X16 iovss sg13g2_Clamp_N43N43D4R_0.gate.t43 iovdd.t29 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X17 iovdd.t109 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t19 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X18 iovdd.t117 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t18 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X19 iovss sg13g2_Clamp_N43N43D4R_0.gate.t44 iovdd.t69 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X20 iovdd.t60 sg13g2_Clamp_N43N43D4R_0.gate.t45 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X21 iovss sg13g2_Clamp_N43N43D4R_0.gate.t46 iovdd.t26 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X22 iovss sg13g2_Clamp_N43N43D4R_0.gate.t47 iovdd.t84 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X23 iovss sg13g2_Clamp_N43N43D4R_0.gate.t48 iovdd.t23 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X24 iovdd.t58 sg13g2_Clamp_N43N43D4R_0.gate.t49 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X25 sg13g2_Clamp_N43N43D4R_0.gate.t3 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t108 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X26 a_11365_11542# a_11695_7456# iovss rppd l=20u w=1u
X27 iovdd.t113 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t20 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X28 iovss sg13g2_Clamp_N43N43D4R_0.gate.t50 iovdd.t19 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X29 sg13g2_Clamp_N43N43D4R_0.gate.t8 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t91 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X30 a_8725_11542# a_9055_7456# iovss rppd l=20u w=1u
X31 iovdd.t79 sg13g2_Clamp_N43N43D4R_0.gate.t51 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X32 iovdd.t78 sg13g2_Clamp_N43N43D4R_0.gate.t52 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X33 iovss sg13g2_Clamp_N43N43D4R_0.gate.t53 iovdd.t54 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X34 a_10045_11542# a_9715_7456# iovss rppd l=20u w=1u
X35 iovdd.t53 sg13g2_Clamp_N43N43D4R_0.gate.t54 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X36 iovss sg13g2_Clamp_N43N43D4R_0.gate.t55 iovdd.t82 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X37 iovss sg13g2_Clamp_N43N43D4R_0.gate.t56 iovdd.t52 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X38 iovdd.t50 sg13g2_Clamp_N43N43D4R_0.gate.t57 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X39 iovdd.t0 sg13g2_Clamp_N43N43D4R_0.gate.t58 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X40 iovss sg13g2_Clamp_N43N43D4R_0.gate.t59 iovdd.t14 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X41 iovdd.t122 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t23 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X42 iovss sg13g2_Clamp_N43N43D4R_0.gate.t60 iovdd.t12 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X43 sg13g2_Clamp_N43N43D4R_0.gate.t14 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t131 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X44 iovss sg13g2_RCClampResistor_0.pin2.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=2.24759n ps=2.5228m w=9u l=9.5u
X45 iovss sg13g2_Clamp_N43N43D4R_0.gate.t61 iovdd.t9 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X46 iovss sg13g2_RCClampResistor_0.pin2.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X47 iovss sg13g2_Clamp_N43N43D4R_0.gate.t62 iovdd.t45 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X48 a_4105_11542# a_4435_7456# iovss rppd l=20u w=1u
X49 a_7405_11542# a_7735_7456# iovss rppd l=20u w=1u
X50 iovdd.t73 sg13g2_Clamp_N43N43D4R_0.gate.t63 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X51 iovdd.t31 sg13g2_Clamp_N43N43D4R_0.gate.t64 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X52 iovss sg13g2_Clamp_N43N43D4R_0.gate.t31 iovdd.t44 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X53 iovdd.t86 sg13g2_Clamp_N43N43D4R_0.gate.t65 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X54 iovdd.t85 sg13g2_Clamp_N43N43D4R_0.gate.t66 iovss iovss sg13_hv_nmos ad=3.256p pd=10.28u as=1.408p ps=5.04u w=4.4u l=0.6u
X55 iovss sg13g2_Clamp_N43N43D4R_0.gate.t34 iovdd.t1 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X56 iovdd.t72 sg13g2_Clamp_N43N43D4R_0.gate.t67 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X57 iovdd.t71 sg13g2_Clamp_N43N43D4R_0.gate.t68 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X58 sg13g2_Clamp_N43N43D4R_0.gate.t22 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t97 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X59 sg13g2_Clamp_N43N43D4R_0.gate.t16 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t104 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X60 iovss sg13g2_Clamp_N43N43D4R_0.gate.t69 iovdd.t41 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X61 iovss sg13g2_RCClampResistor_0.pin2.t2 sg13g2_Clamp_N43N43D4R_0.gate.t28 iovss sg13_hv_nmos ad=1.71p pd=9.38u as=1.71p ps=9.38u w=9u l=0.5u
X62 iovss sg13g2_Clamp_N43N43D4R_0.gate.t70 iovdd.t13 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X63 iovss sg13g2_Clamp_N43N43D4R_0.gate.t71 iovdd.t51 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X64 iovdd.t84 sg13g2_Clamp_N43N43D4R_0.gate.t72 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X65 sg13g2_Clamp_N43N43D4R_0.gate.t11 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t103 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X66 iovss sg13g2_RCClampResistor_0.pin2.t2 sg13g2_Clamp_N43N43D4R_0.gate.t27 iovss sg13_hv_nmos ad=1.71p pd=9.38u as=1.71p ps=9.38u w=9u l=0.5u
X67 sg13g2_Clamp_N43N43D4R_0.gate.t9 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t102 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X68 iovss sg13g2_RCClampResistor_0.pin2.t2 sg13g2_Clamp_N43N43D4R_0.gate.t26 iovss sg13_hv_nmos ad=1.71p pd=9.38u as=1.71p ps=9.38u w=9u l=0.5u
X69 iovss sg13g2_RCClampResistor_0.pin2.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X70 iovss sg13g2_Clamp_N43N43D4R_0.gate.t73 iovdd.t83 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X71 iovdd.t67 sg13g2_Clamp_N43N43D4R_0.gate.t74 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X72 iovdd.t65 sg13g2_Clamp_N43N43D4R_0.gate.t75 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X73 sg13g2_Clamp_N43N43D4R_0.gate.t7 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t101 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X74 iovss sg13g2_RCClampResistor_0.pin2.t2 sg13g2_Clamp_N43N43D4R_0.gate.t25 iovss sg13_hv_nmos ad=1.71p pd=9.38u as=1.71p ps=9.38u w=9u l=0.5u
X75 iovss sg13g2_RCClampResistor_0.pin2.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X76 iovdd.t83 sg13g2_Clamp_N43N43D4R_0.gate.t76 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=2.068p ps=9.74u w=4.4u l=0.6u
X77 sg13g2_Clamp_N43N43D4R_0.gate.t12 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t100 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X78 iovss sg13g2_RCClampResistor_0.pin2.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X79 iovdd.t64 sg13g2_Clamp_N43N43D4R_0.gate.t77 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X80 iovss sg13g2_Clamp_N43N43D4R_0.gate.t78 iovdd.t32 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X81 a_4765_11542# a_5095_7456# iovss rppd l=20u w=1u
X82 a_8065_11542# a_8395_7456# iovss rppd l=20u w=1u
X83 iovdd.t36 sg13g2_Clamp_N43N43D4R_0.gate.t45 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X84 iovdd.t18 sg13g2_Clamp_N43N43D4R_0.gate.t79 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X85 iovdd.t63 sg13g2_Clamp_N43N43D4R_0.gate.t80 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X86 iovss sg13g2_RCClampResistor_0.pin2.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X87 iovdd.t15 sg13g2_Clamp_N43N43D4R_0.gate.t81 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X88 sg13g2_Clamp_N43N43D4R_0.gate.t5 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t111 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X89 iovdd.t82 sg13g2_Clamp_N43N43D4R_0.gate.t82 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X90 sg13g2_Clamp_N43N43D4R_0.gate.t15 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t106 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X91 iovss sg13g2_Clamp_N43N43D4R_0.gate.t83 iovdd.t81 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X92 sg13g2_Clamp_N43N43D4R_0.gate.t19 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t122 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X93 iovss sg13g2_RCClampResistor_0.pin2.t2 sg13g2_Clamp_N43N43D4R_0.gate.t30 iovss sg13_hv_nmos ad=1.71p pd=9.38u as=1.71p ps=9.38u w=9u l=0.5u
X94 iovdd.t81 sg13g2_Clamp_N43N43D4R_0.gate.t84 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X95 iovss sg13g2_Clamp_N43N43D4R_0.gate.t85 iovdd.t80 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X96 iovdd.t61 sg13g2_Clamp_N43N43D4R_0.gate.t86 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X97 sg13g2_Clamp_N43N43D4R_0.gate.t0 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t105 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X98 sg13g2_Clamp_N43N43D4R_0.gate.t1 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t96 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X99 iovss sg13g2_RCClampResistor_0.pin2.t2 sg13g2_Clamp_N43N43D4R_0.gate.t29 iovss sg13_hv_nmos ad=1.71p pd=9.38u as=1.71p ps=9.38u w=9u l=0.5u
X100 iovdd.t59 sg13g2_Clamp_N43N43D4R_0.gate.t52 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X101 iovdd.t10 sg13g2_Clamp_N43N43D4R_0.gate.t87 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X102 iovdd.t25 sg13g2_Clamp_N43N43D4R_0.gate.t54 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X103 a_10705_11542# a_11035_7456# iovss rppd l=20u w=1u
X104 iovdd.t46 sg13g2_Clamp_N43N43D4R_0.gate.t88 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X105 sg13g2_Clamp_N43N43D4R_0.gate.t6 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t94 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X106 iovdd.t57 sg13g2_Clamp_N43N43D4R_0.gate.t89 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X107 sg13g2_Clamp_N43N43D4R_0.gate.t17 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t90 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X108 iovdd.t88 a_3775_7456# iovss rppd l=20u w=1u
X109 iovss sg13g2_Clamp_N43N43D4R_0.gate.t90 iovdd.t34 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X110 sg13g2_Clamp_N43N43D4R_0.gate.t24 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t117 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X111 iovss sg13g2_Clamp_N43N43D4R_0.gate.t37 iovdd.t79 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X112 iovss sg13g2_Clamp_N43N43D4R_0.gate.t91 iovdd.t78 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X113 sg13g2_Clamp_N43N43D4R_0.gate.t4 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t92 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X114 iovss sg13g2_Clamp_N43N43D4R_0.gate.t92 iovdd.t77 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X115 sg13g2_Clamp_N43N43D4R_0.gate.t23 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t115 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X116 iovdd.t77 sg13g2_Clamp_N43N43D4R_0.gate.t93 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X117 iovss sg13g2_Clamp_N43N43D4R_0.gate.t94 iovdd.t75 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X118 a_5425_11542# a_5095_7456# iovss rppd l=20u w=1u
X119 a_8725_11542# a_8395_7456# iovss rppd l=20u w=1u
X120 iovdd.t76 sg13g2_Clamp_N43N43D4R_0.gate.t66 iovss iovss sg13_hv_nmos ad=3.256p pd=10.28u as=1.408p ps=5.04u w=4.4u l=0.6u
X121 iovdd.t75 sg13g2_Clamp_N43N43D4R_0.gate.t95 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X122 iovdd.t47 sg13g2_Clamp_N43N43D4R_0.gate.t96 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X123 iovdd.t48 sg13g2_Clamp_N43N43D4R_0.gate.t67 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X124 iovdd.t74 sg13g2_Clamp_N43N43D4R_0.gate.t97 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X125 iovss sg13g2_Clamp_N43N43D4R_0.gate.t44 iovdd.t24 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X126 iovss sg13g2_Clamp_N43N43D4R_0.gate.t48 iovdd.t73 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X127 iovss sg13g2_Clamp_N43N43D4R_0.gate.t98 iovdd.t56 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X128 iovss sg13g2_Clamp_N43N43D4R_0.gate.t71 iovdd.t21 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X129 iovdd.t6 sg13g2_Clamp_N43N43D4R_0.gate.t33 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X130 sg13g2_Clamp_N43N43D4R_0.gate.t10 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t114 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=2.38p ps=14.68u w=7u l=0.5u
X131 iovss sg13g2_RCClampResistor_0.pin2.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X132 iovss sg13g2_RCClampResistor_0.pin2.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X133 iovss sg13g2_Clamp_N43N43D4R_0.gate.t36 iovdd.t72 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X134 iovss sg13g2_Clamp_N43N43D4R_0.gate.t73 iovdd.t70 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X135 iovdd.t43 sg13g2_Clamp_N43N43D4R_0.gate.t74 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X136 iovss sg13g2_Clamp_N43N43D4R_0.gate.t99 iovdd.t71 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X137 iovdd.t70 sg13g2_Clamp_N43N43D4R_0.gate.t76 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=2.068p ps=9.74u w=4.4u l=0.6u
X138 iovdd.t42 sg13g2_Clamp_N43N43D4R_0.gate.t77 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X139 iovdd.t69 sg13g2_Clamp_N43N43D4R_0.gate.t79 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X140 a_6085_11542# a_5755_7456# iovss rppd l=20u w=1u
X141 a_9385_11542# a_9055_7456# iovss rppd l=20u w=1u
X142 iovss sg13g2_Clamp_N43N43D4R_0.gate.t41 iovdd.t49 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X143 iovss sg13g2_Clamp_N43N43D4R_0.gate.t56 iovdd.t68 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X144 iovss sg13g2_Clamp_N43N43D4R_0.gate.t43 iovdd.t67 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X145 iovdd.t66 sg13g2_Clamp_N43N43D4R_0.gate.t42 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X146 iovss sg13g2_Clamp_N43N43D4R_0.gate.t60 iovdd.t65 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X147 a_10045_11542# a_10375_7456# iovss rppd l=20u w=1u
X148 sg13g2_Clamp_N43N43D4R_0.gate.t21 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t113 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X149 iovss sg13g2_Clamp_N43N43D4R_0.gate.t46 iovdd.t64 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X150 iovss sg13g2_Clamp_N43N43D4R_0.gate.t100 iovdd.t8 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X151 sg13g2_Clamp_N43N43D4R_0.gate.t13 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t99 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X152 iovss sg13g2_Clamp_N43N43D4R_0.gate.t101 iovdd.t63 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X153 iovdd.t111 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t4 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X154 sg13g2_Clamp_N43N43D4R_0.gate.t2 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t98 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X155 iovdd.t17 sg13g2_Clamp_N43N43D4R_0.gate.t88 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X156 iovss sg13g2_Clamp_N43N43D4R_0.gate.t31 iovdd.t62 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X157 sg13g2_RCClampResistor_0.pin2.t0 a_11695_7456# iovss rppd l=20u w=1u
X158 iovss sg13g2_Clamp_N43N43D4R_0.gate.t90 iovdd.t2 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X159 iovss sg13g2_Clamp_N43N43D4R_0.gate.t34 iovdd.t61 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X160 iovdd.t28 sg13g2_Clamp_N43N43D4R_0.gate.t51 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X161 sg13g2_Clamp_N43N43D4R_0.gate.t18 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t109 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X162 a_4765_11542# a_4435_7456# iovss rppd l=20u w=1u
X163 iovss sg13g2_Clamp_N43N43D4R_0.gate.t53 iovdd.t60 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X164 iovss sg13g2_Clamp_N43N43D4R_0.gate.t91 iovdd.t59 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X165 iovss sg13g2_Clamp_N43N43D4R_0.gate.t102 iovdd.t58 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X166 iovdd.t108 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t2 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X167 iovss sg13g2_Clamp_N43N43D4R_0.gate.t92 iovdd.t55 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X168 iovss sg13g2_Clamp_N43N43D4R_0.gate.t103 iovdd.t57 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X169 iovdd.t56 sg13g2_Clamp_N43N43D4R_0.gate.t58 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X170 sg13g2_Clamp_N43N43D4R_0.gate.t20 sg13g2_RCClampResistor_0.pin2.t1 iovdd.t95 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X171 iovdd.t55 sg13g2_Clamp_N43N43D4R_0.gate.t93 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X172 a_9385_11542# a_9715_7456# iovss rppd l=20u w=1u
X173 iovss sg13g2_RCClampResistor_0.pin2.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X174 a_6085_11542# a_6415_7456# iovss rppd l=20u w=1u
X175 iovdd.t54 sg13g2_Clamp_N43N43D4R_0.gate.t45 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X176 iovss sg13g2_RCClampResistor_0.pin2.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X177 a_10705_11542# a_10375_7456# iovss rppd l=20u w=1u
X178 iovss sg13g2_Clamp_N43N43D4R_0.gate.t98 iovdd.t30 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X179 iovss sg13g2_Clamp_N43N43D4R_0.gate.t62 iovdd.t53 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X180 iovdd.t52 sg13g2_Clamp_N43N43D4R_0.gate.t33 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X181 iovdd.t51 sg13g2_Clamp_N43N43D4R_0.gate.t64 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X182 iovdd.t16 sg13g2_Clamp_N43N43D4R_0.gate.t63 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X183 iovss sg13g2_Clamp_N43N43D4R_0.gate.t104 iovdd.t50 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X184 iovdd.t49 sg13g2_Clamp_N43N43D4R_0.gate.t65 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X185 iovss sg13g2_Clamp_N43N43D4R_0.gate.t36 iovdd.t48 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X186 iovss sg13g2_Clamp_N43N43D4R_0.gate.t105 iovdd.t47 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X187 iovdd.t106 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t14 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X188 iovss sg13g2_Clamp_N43N43D4R_0.gate.t70 iovdd.t46 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X189 iovdd.t7 sg13g2_Clamp_N43N43D4R_0.gate.t52 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X190 iovdd.t105 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t13 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X191 iovdd.t45 sg13g2_Clamp_N43N43D4R_0.gate.t54 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X192 iovss sg13g2_Clamp_N43N43D4R_0.gate.t41 iovdd.t20 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X193 a_6745_11542# a_7075_7456# iovss rppd l=20u w=1u
X194 iovdd.t44 sg13g2_Clamp_N43N43D4R_0.gate.t42 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X195 iovss sg13g2_Clamp_N43N43D4R_0.gate.t43 iovdd.t43 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X196 iovdd.t5 sg13g2_Clamp_N43N43D4R_0.gate.t75 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X197 iovdd.t104 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t22 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X198 a_11365_11542# a_11035_7456# iovss rppd l=20u w=1u
X199 iovss sg13g2_Clamp_N43N43D4R_0.gate.t46 iovdd.t42 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X200 iovdd.t41 sg13g2_Clamp_N43N43D4R_0.gate.t106 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X201 sg13g2_Clamp_N43N43D4R_0.gate.t28 sg13g2_RCClampResistor_0.pin2.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=1.71p ps=9.38u w=9u l=0.5u
X202 iovss sg13g2_RCClampResistor_0.pin2.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X203 iovdd.t103 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t1 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X204 sg13g2_Clamp_N43N43D4R_0.gate.t27 sg13g2_RCClampResistor_0.pin2.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=1.71p ps=9.38u w=9u l=0.5u
X205 iovss sg13g2_RCClampResistor_0.pin2.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X206 iovdd.t102 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t8 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X207 sg13g2_Clamp_N43N43D4R_0.gate.t26 sg13g2_RCClampResistor_0.pin2.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=3.06p ps=18.68u w=9u l=0.5u
X208 iovss sg13g2_Clamp_N43N43D4R_0.gate.t83 iovdd.t40 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X209 sg13g2_Clamp_N43N43D4R_0.gate.t25 sg13g2_RCClampResistor_0.pin2.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=3.06p ps=18.68u w=9u l=0.5u
X210 iovdd.t40 sg13g2_Clamp_N43N43D4R_0.gate.t84 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X211 iovdd.t39 sg13g2_Clamp_N43N43D4R_0.gate.t66 iovss iovss sg13_hv_nmos ad=3.256p pd=10.28u as=1.408p ps=5.04u w=4.4u l=0.6u
X212 iovdd.t101 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t6 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X213 iovdd.t38 sg13g2_Clamp_N43N43D4R_0.gate.t86 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X214 iovdd.t37 sg13g2_Clamp_N43N43D4R_0.gate.t67 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X215 iovdd.t100 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t17 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X216 iovdd.t99 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t12 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X217 iovss sg13g2_Clamp_N43N43D4R_0.gate.t53 iovdd.t36 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X218 iovdd.t35 sg13g2_Clamp_N43N43D4R_0.gate.t51 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X219 iovdd.t34 sg13g2_Clamp_N43N43D4R_0.gate.t87 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X220 iovdd.t33 sg13g2_Clamp_N43N43D4R_0.gate.t107 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X221 a_5425_11542# a_5755_7456# iovss rppd l=20u w=1u
X222 iovdd.t32 sg13g2_Clamp_N43N43D4R_0.gate.t108 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X223 iovss sg13g2_Clamp_N43N43D4R_0.gate.t71 iovdd.t31 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X224 iovdd.t98 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t5 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X225 iovdd.t30 sg13g2_Clamp_N43N43D4R_0.gate.t58 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X226 iovdd.t97 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t15 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X227 iovss sg13g2_RCClampResistor_0.pin2.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X228 iovdd.t29 sg13g2_Clamp_N43N43D4R_0.gate.t74 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X229 iovss sg13g2_Clamp_N43N43D4R_0.gate.t73 iovdd.t27 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X230 iovss sg13g2_Clamp_N43N43D4R_0.gate.t37 iovdd.t28 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X231 iovss sg13g2_RCClampResistor_0.pin2.t2 iovss iovss sg13_hv_nmos ad=1.71p pd=9.38u as=0 ps=0 w=9u l=9.5u
X232 a_4105_11542# a_3775_7456# iovss rppd l=20u w=1u
X233 a_7405_11542# a_7075_7456# iovss rppd l=20u w=1u
X234 iovdd.t27 sg13g2_Clamp_N43N43D4R_0.gate.t76 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=2.068p ps=9.74u w=4.4u l=0.6u
X235 iovdd.t96 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t0 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X236 iovdd.t26 sg13g2_Clamp_N43N43D4R_0.gate.t77 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X237 iovss sg13g2_Clamp_N43N43D4R_0.gate.t62 iovdd.t25 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X238 iovdd.t24 sg13g2_Clamp_N43N43D4R_0.gate.t79 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X239 iovdd.t95 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t7 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X240 iovdd.t23 sg13g2_Clamp_N43N43D4R_0.gate.t63 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X241 iovdd.t22 sg13g2_Clamp_N43N43D4R_0.gate.t109 iovss iovss sg13_hv_nmos ad=3.256p pd=10.28u as=1.408p ps=5.04u w=4.4u l=0.6u
X242 iovdd.t94 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t3 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X243 iovdd.t21 sg13g2_Clamp_N43N43D4R_0.gate.t64 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X244 iovdd.t20 sg13g2_Clamp_N43N43D4R_0.gate.t65 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X245 iovdd.t19 sg13g2_Clamp_N43N43D4R_0.gate.t110 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X246 iovdd.t93 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t24 iovdd.t89 sg13_hv_pmos ad=2.38p pd=14.68u as=1.33p ps=7.38u w=7u l=0.5u
X247 iovss sg13g2_Clamp_N43N43D4R_0.gate.t44 iovdd.t18 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X248 iovss sg13g2_Clamp_N43N43D4R_0.gate.t70 iovdd.t17 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X249 iovss sg13g2_Clamp_N43N43D4R_0.gate.t48 iovdd.t16 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X250 iovss sg13g2_Clamp_N43N43D4R_0.gate.t111 iovdd.t15 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X251 iovdd.t92 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t11 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X252 iovdd.t14 sg13g2_Clamp_N43N43D4R_0.gate.t112 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X253 iovdd.t13 sg13g2_Clamp_N43N43D4R_0.gate.t88 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X254 a_8065_11542# a_7735_7456# iovss rppd l=20u w=1u
X255 iovss sg13g2_Clamp_N43N43D4R_0.gate.t113 iovdd.t11 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X256 iovdd.t12 sg13g2_Clamp_N43N43D4R_0.gate.t75 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X257 iovdd.t11 sg13g2_Clamp_N43N43D4R_0.gate.t114 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=2.068p ps=9.74u w=4.4u l=0.6u
X258 iovss sg13g2_Clamp_N43N43D4R_0.gate.t90 iovdd.t10 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X259 iovdd.t9 sg13g2_Clamp_N43N43D4R_0.gate.t115 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X260 iovdd.t8 sg13g2_Clamp_N43N43D4R_0.gate.t116 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X261 iovss sg13g2_Clamp_N43N43D4R_0.gate.t91 iovdd.t7 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X262 iovss sg13g2_Clamp_N43N43D4R_0.gate.t117 dantenna l=0.48u w=0.48u
X263 iovss sg13g2_Clamp_N43N43D4R_0.gate.t56 iovdd.t6 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X264 iovss sg13g2_Clamp_N43N43D4R_0.gate.t92 iovdd.t4 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X265 iovdd.t91 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t10 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X266 iovss sg13g2_Clamp_N43N43D4R_0.gate.t60 iovdd.t5 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X267 iovss sg13g2_Clamp_N43N43D4R_0.gate.t83 iovdd.t3 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X268 iovdd.t4 sg13g2_Clamp_N43N43D4R_0.gate.t93 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X269 iovdd.t90 sg13g2_RCClampResistor_0.pin2.t1 sg13g2_Clamp_N43N43D4R_0.gate.t16 iovdd.t89 sg13_hv_pmos ad=1.33p pd=7.38u as=1.33p ps=7.38u w=7u l=0.5u
X270 iovdd.t3 sg13g2_Clamp_N43N43D4R_0.gate.t84 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X271 iovdd.t2 sg13g2_Clamp_N43N43D4R_0.gate.t87 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X272 iovdd.t1 sg13g2_Clamp_N43N43D4R_0.gate.t86 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X273 a_6745_11542# a_6415_7456# iovss rppd l=20u w=1u
X274 iovss sg13g2_Clamp_N43N43D4R_0.gate.t98 iovdd.t0 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
R0 sg13g2_Clamp_N43N43D4R_0.gate.n85 sg13g2_Clamp_N43N43D4R_0.gate.t117 17.2912
R1 sg13g2_Clamp_N43N43D4R_0.gate.n2 sg13g2_Clamp_N43N43D4R_0.gate.n0 6.58671
R2 sg13g2_Clamp_N43N43D4R_0.gate.n82 sg13g2_Clamp_N43N43D4R_0.gate.n81 5.73421
R3 sg13g2_Clamp_N43N43D4R_0.gate.n80 sg13g2_Clamp_N43N43D4R_0.gate.n79 5.73421
R4 sg13g2_Clamp_N43N43D4R_0.gate.n78 sg13g2_Clamp_N43N43D4R_0.gate.n77 5.73421
R5 sg13g2_Clamp_N43N43D4R_0.gate.n76 sg13g2_Clamp_N43N43D4R_0.gate.n75 5.73421
R6 sg13g2_Clamp_N43N43D4R_0.gate.n74 sg13g2_Clamp_N43N43D4R_0.gate.n73 5.73421
R7 sg13g2_Clamp_N43N43D4R_0.gate.n72 sg13g2_Clamp_N43N43D4R_0.gate.n71 5.73421
R8 sg13g2_Clamp_N43N43D4R_0.gate.n70 sg13g2_Clamp_N43N43D4R_0.gate.n69 5.73421
R9 sg13g2_Clamp_N43N43D4R_0.gate.n68 sg13g2_Clamp_N43N43D4R_0.gate.n67 5.73421
R10 sg13g2_Clamp_N43N43D4R_0.gate.n66 sg13g2_Clamp_N43N43D4R_0.gate.n65 5.73421
R11 sg13g2_Clamp_N43N43D4R_0.gate.n64 sg13g2_Clamp_N43N43D4R_0.gate.n63 5.73421
R12 sg13g2_Clamp_N43N43D4R_0.gate.n62 sg13g2_Clamp_N43N43D4R_0.gate.n61 5.73421
R13 sg13g2_Clamp_N43N43D4R_0.gate.n60 sg13g2_Clamp_N43N43D4R_0.gate.n59 5.73421
R14 sg13g2_Clamp_N43N43D4R_0.gate.n58 sg13g2_Clamp_N43N43D4R_0.gate.n57 5.73421
R15 sg13g2_Clamp_N43N43D4R_0.gate.n56 sg13g2_Clamp_N43N43D4R_0.gate.n55 5.73421
R16 sg13g2_Clamp_N43N43D4R_0.gate.n54 sg13g2_Clamp_N43N43D4R_0.gate.n53 5.73421
R17 sg13g2_Clamp_N43N43D4R_0.gate.n52 sg13g2_Clamp_N43N43D4R_0.gate.n51 5.73421
R18 sg13g2_Clamp_N43N43D4R_0.gate.n50 sg13g2_Clamp_N43N43D4R_0.gate.n49 5.73421
R19 sg13g2_Clamp_N43N43D4R_0.gate.n48 sg13g2_Clamp_N43N43D4R_0.gate.n47 5.73421
R20 sg13g2_Clamp_N43N43D4R_0.gate.n46 sg13g2_Clamp_N43N43D4R_0.gate.n45 5.73421
R21 sg13g2_Clamp_N43N43D4R_0.gate.n44 sg13g2_Clamp_N43N43D4R_0.gate.n43 5.73421
R22 sg13g2_Clamp_N43N43D4R_0.gate.n42 sg13g2_Clamp_N43N43D4R_0.gate.n41 5.73421
R23 sg13g2_Clamp_N43N43D4R_0.gate.n40 sg13g2_Clamp_N43N43D4R_0.gate.n39 5.73421
R24 sg13g2_Clamp_N43N43D4R_0.gate.n38 sg13g2_Clamp_N43N43D4R_0.gate.n37 5.73421
R25 sg13g2_Clamp_N43N43D4R_0.gate.n36 sg13g2_Clamp_N43N43D4R_0.gate.n35 5.73421
R26 sg13g2_Clamp_N43N43D4R_0.gate.n34 sg13g2_Clamp_N43N43D4R_0.gate.n33 5.73421
R27 sg13g2_Clamp_N43N43D4R_0.gate.n32 sg13g2_Clamp_N43N43D4R_0.gate.n31 5.73421
R28 sg13g2_Clamp_N43N43D4R_0.gate.n30 sg13g2_Clamp_N43N43D4R_0.gate.n29 5.73421
R29 sg13g2_Clamp_N43N43D4R_0.gate.n28 sg13g2_Clamp_N43N43D4R_0.gate.n27 5.73421
R30 sg13g2_Clamp_N43N43D4R_0.gate.n26 sg13g2_Clamp_N43N43D4R_0.gate.n25 5.73421
R31 sg13g2_Clamp_N43N43D4R_0.gate.n24 sg13g2_Clamp_N43N43D4R_0.gate.n23 5.73421
R32 sg13g2_Clamp_N43N43D4R_0.gate.n22 sg13g2_Clamp_N43N43D4R_0.gate.n21 5.73421
R33 sg13g2_Clamp_N43N43D4R_0.gate.n20 sg13g2_Clamp_N43N43D4R_0.gate.n19 5.73421
R34 sg13g2_Clamp_N43N43D4R_0.gate.n18 sg13g2_Clamp_N43N43D4R_0.gate.n17 5.73421
R35 sg13g2_Clamp_N43N43D4R_0.gate.n16 sg13g2_Clamp_N43N43D4R_0.gate.n15 5.73421
R36 sg13g2_Clamp_N43N43D4R_0.gate.n14 sg13g2_Clamp_N43N43D4R_0.gate.n13 5.73421
R37 sg13g2_Clamp_N43N43D4R_0.gate.n12 sg13g2_Clamp_N43N43D4R_0.gate.n11 5.73421
R38 sg13g2_Clamp_N43N43D4R_0.gate.n10 sg13g2_Clamp_N43N43D4R_0.gate.n9 5.73421
R39 sg13g2_Clamp_N43N43D4R_0.gate.n8 sg13g2_Clamp_N43N43D4R_0.gate.n7 5.73421
R40 sg13g2_Clamp_N43N43D4R_0.gate.n6 sg13g2_Clamp_N43N43D4R_0.gate.n5 5.73421
R41 sg13g2_Clamp_N43N43D4R_0.gate.n4 sg13g2_Clamp_N43N43D4R_0.gate.n3 5.73421
R42 sg13g2_Clamp_N43N43D4R_0.gate.n2 sg13g2_Clamp_N43N43D4R_0.gate.n1 5.73421
R43 sg13g2_Clamp_N43N43D4R_0.gate.n84 sg13g2_Clamp_N43N43D4R_0.gate.n83 5.73421
R44 sg13g2_Clamp_N43N43D4R_0.gate sg13g2_Clamp_N43N43D4R_0.gate.n85 4.50322
R45 sg13g2_Clamp_N43N43D4R_0.gate.n85 sg13g2_Clamp_N43N43D4R_0.gate.n84 2.48679
R46 sg13g2_Clamp_N43N43D4R_0.gate.n86 sg13g2_Clamp_N43N43D4R_0.gate.t24 1.72119
R47 sg13g2_Clamp_N43N43D4R_0.gate.n98 sg13g2_Clamp_N43N43D4R_0.gate.t1 1.70127
R48 sg13g2_Clamp_N43N43D4R_0.gate.n108 sg13g2_Clamp_N43N43D4R_0.gate.t8 1.69835
R49 sg13g2_Clamp_N43N43D4R_0.gate.n107 sg13g2_Clamp_N43N43D4R_0.gate.t9 1.69835
R50 sg13g2_Clamp_N43N43D4R_0.gate.n106 sg13g2_Clamp_N43N43D4R_0.gate.t14 1.69835
R51 sg13g2_Clamp_N43N43D4R_0.gate.n105 sg13g2_Clamp_N43N43D4R_0.gate.t15 1.69835
R52 sg13g2_Clamp_N43N43D4R_0.gate.n104 sg13g2_Clamp_N43N43D4R_0.gate.t22 1.69835
R53 sg13g2_Clamp_N43N43D4R_0.gate.n103 sg13g2_Clamp_N43N43D4R_0.gate.t16 1.69835
R54 sg13g2_Clamp_N43N43D4R_0.gate.n102 sg13g2_Clamp_N43N43D4R_0.gate.t17 1.69835
R55 sg13g2_Clamp_N43N43D4R_0.gate.n101 sg13g2_Clamp_N43N43D4R_0.gate.t12 1.69835
R56 sg13g2_Clamp_N43N43D4R_0.gate.n100 sg13g2_Clamp_N43N43D4R_0.gate.t13 1.69835
R57 sg13g2_Clamp_N43N43D4R_0.gate.n99 sg13g2_Clamp_N43N43D4R_0.gate.t0 1.69835
R58 sg13g2_Clamp_N43N43D4R_0.gate.n97 sg13g2_Clamp_N43N43D4R_0.gate.t11 1.69835
R59 sg13g2_Clamp_N43N43D4R_0.gate.n96 sg13g2_Clamp_N43N43D4R_0.gate.t4 1.69835
R60 sg13g2_Clamp_N43N43D4R_0.gate.n95 sg13g2_Clamp_N43N43D4R_0.gate.t5 1.69835
R61 sg13g2_Clamp_N43N43D4R_0.gate.n94 sg13g2_Clamp_N43N43D4R_0.gate.t2 1.69835
R62 sg13g2_Clamp_N43N43D4R_0.gate.n93 sg13g2_Clamp_N43N43D4R_0.gate.t3 1.69835
R63 sg13g2_Clamp_N43N43D4R_0.gate.n92 sg13g2_Clamp_N43N43D4R_0.gate.t6 1.69835
R64 sg13g2_Clamp_N43N43D4R_0.gate.n91 sg13g2_Clamp_N43N43D4R_0.gate.t7 1.69835
R65 sg13g2_Clamp_N43N43D4R_0.gate.n90 sg13g2_Clamp_N43N43D4R_0.gate.t20 1.69835
R66 sg13g2_Clamp_N43N43D4R_0.gate.n89 sg13g2_Clamp_N43N43D4R_0.gate.t21 1.69835
R67 sg13g2_Clamp_N43N43D4R_0.gate.n88 sg13g2_Clamp_N43N43D4R_0.gate.t23 1.69835
R68 sg13g2_Clamp_N43N43D4R_0.gate.n87 sg13g2_Clamp_N43N43D4R_0.gate.t19 1.69835
R69 sg13g2_Clamp_N43N43D4R_0.gate.n86 sg13g2_Clamp_N43N43D4R_0.gate.t18 1.69835
R70 sg13g2_Clamp_N43N43D4R_0.gate.n109 sg13g2_Clamp_N43N43D4R_0.gate.t10 1.69585
R71 sg13g2_Clamp_N43N43D4R_0.gate.n110 sg13g2_Clamp_N43N43D4R_0.gate.t25 1.43866
R72 sg13g2_Clamp_N43N43D4R_0.gate.n110 sg13g2_Clamp_N43N43D4R_0.gate.t29 1.43866
R73 sg13g2_Clamp_N43N43D4R_0.gate.n110 sg13g2_Clamp_N43N43D4R_0.gate.t27 1.43866
R74 sg13g2_Clamp_N43N43D4R_0.gate.n111 sg13g2_Clamp_N43N43D4R_0.gate.t26 1.43866
R75 sg13g2_Clamp_N43N43D4R_0.gate.n111 sg13g2_Clamp_N43N43D4R_0.gate.t30 1.43866
R76 sg13g2_Clamp_N43N43D4R_0.gate.n111 sg13g2_Clamp_N43N43D4R_0.gate.t28 1.43866
R77 sg13g2_Clamp_N43N43D4R_0.gate.n4 sg13g2_Clamp_N43N43D4R_0.gate.n2 1.22425
R78 sg13g2_Clamp_N43N43D4R_0.gate.n8 sg13g2_Clamp_N43N43D4R_0.gate.n6 1.22425
R79 sg13g2_Clamp_N43N43D4R_0.gate.n12 sg13g2_Clamp_N43N43D4R_0.gate.n10 1.22425
R80 sg13g2_Clamp_N43N43D4R_0.gate.n16 sg13g2_Clamp_N43N43D4R_0.gate.n14 1.22425
R81 sg13g2_Clamp_N43N43D4R_0.gate.n20 sg13g2_Clamp_N43N43D4R_0.gate.n18 1.22425
R82 sg13g2_Clamp_N43N43D4R_0.gate.n24 sg13g2_Clamp_N43N43D4R_0.gate.n22 1.22425
R83 sg13g2_Clamp_N43N43D4R_0.gate.n28 sg13g2_Clamp_N43N43D4R_0.gate.n26 1.22425
R84 sg13g2_Clamp_N43N43D4R_0.gate.n32 sg13g2_Clamp_N43N43D4R_0.gate.n30 1.22425
R85 sg13g2_Clamp_N43N43D4R_0.gate.n36 sg13g2_Clamp_N43N43D4R_0.gate.n34 1.22425
R86 sg13g2_Clamp_N43N43D4R_0.gate.n40 sg13g2_Clamp_N43N43D4R_0.gate.n38 1.22425
R87 sg13g2_Clamp_N43N43D4R_0.gate.n44 sg13g2_Clamp_N43N43D4R_0.gate.n42 1.22425
R88 sg13g2_Clamp_N43N43D4R_0.gate.n48 sg13g2_Clamp_N43N43D4R_0.gate.n46 1.22425
R89 sg13g2_Clamp_N43N43D4R_0.gate.n52 sg13g2_Clamp_N43N43D4R_0.gate.n50 1.22425
R90 sg13g2_Clamp_N43N43D4R_0.gate.n56 sg13g2_Clamp_N43N43D4R_0.gate.n54 1.22425
R91 sg13g2_Clamp_N43N43D4R_0.gate.n60 sg13g2_Clamp_N43N43D4R_0.gate.n58 1.22425
R92 sg13g2_Clamp_N43N43D4R_0.gate.n64 sg13g2_Clamp_N43N43D4R_0.gate.n62 1.22425
R93 sg13g2_Clamp_N43N43D4R_0.gate.n68 sg13g2_Clamp_N43N43D4R_0.gate.n66 1.22425
R94 sg13g2_Clamp_N43N43D4R_0.gate.n72 sg13g2_Clamp_N43N43D4R_0.gate.n70 1.22425
R95 sg13g2_Clamp_N43N43D4R_0.gate.n76 sg13g2_Clamp_N43N43D4R_0.gate.n74 1.22425
R96 sg13g2_Clamp_N43N43D4R_0.gate.n80 sg13g2_Clamp_N43N43D4R_0.gate.n78 1.22425
R97 sg13g2_Clamp_N43N43D4R_0.gate.n84 sg13g2_Clamp_N43N43D4R_0.gate.n82 1.22425
R98 sg13g2_Clamp_N43N43D4R_0.gate.n6 sg13g2_Clamp_N43N43D4R_0.gate.n4 0.853
R99 sg13g2_Clamp_N43N43D4R_0.gate.n10 sg13g2_Clamp_N43N43D4R_0.gate.n8 0.853
R100 sg13g2_Clamp_N43N43D4R_0.gate.n14 sg13g2_Clamp_N43N43D4R_0.gate.n12 0.853
R101 sg13g2_Clamp_N43N43D4R_0.gate.n18 sg13g2_Clamp_N43N43D4R_0.gate.n16 0.853
R102 sg13g2_Clamp_N43N43D4R_0.gate.n22 sg13g2_Clamp_N43N43D4R_0.gate.n20 0.853
R103 sg13g2_Clamp_N43N43D4R_0.gate.n26 sg13g2_Clamp_N43N43D4R_0.gate.n24 0.853
R104 sg13g2_Clamp_N43N43D4R_0.gate.n30 sg13g2_Clamp_N43N43D4R_0.gate.n28 0.853
R105 sg13g2_Clamp_N43N43D4R_0.gate.n34 sg13g2_Clamp_N43N43D4R_0.gate.n32 0.853
R106 sg13g2_Clamp_N43N43D4R_0.gate.n38 sg13g2_Clamp_N43N43D4R_0.gate.n36 0.853
R107 sg13g2_Clamp_N43N43D4R_0.gate.n42 sg13g2_Clamp_N43N43D4R_0.gate.n40 0.853
R108 sg13g2_Clamp_N43N43D4R_0.gate.n46 sg13g2_Clamp_N43N43D4R_0.gate.n44 0.853
R109 sg13g2_Clamp_N43N43D4R_0.gate.n50 sg13g2_Clamp_N43N43D4R_0.gate.n48 0.853
R110 sg13g2_Clamp_N43N43D4R_0.gate.n54 sg13g2_Clamp_N43N43D4R_0.gate.n52 0.853
R111 sg13g2_Clamp_N43N43D4R_0.gate.n58 sg13g2_Clamp_N43N43D4R_0.gate.n56 0.853
R112 sg13g2_Clamp_N43N43D4R_0.gate.n62 sg13g2_Clamp_N43N43D4R_0.gate.n60 0.853
R113 sg13g2_Clamp_N43N43D4R_0.gate.n66 sg13g2_Clamp_N43N43D4R_0.gate.n64 0.853
R114 sg13g2_Clamp_N43N43D4R_0.gate.n70 sg13g2_Clamp_N43N43D4R_0.gate.n68 0.853
R115 sg13g2_Clamp_N43N43D4R_0.gate.n74 sg13g2_Clamp_N43N43D4R_0.gate.n72 0.853
R116 sg13g2_Clamp_N43N43D4R_0.gate.n78 sg13g2_Clamp_N43N43D4R_0.gate.n76 0.853
R117 sg13g2_Clamp_N43N43D4R_0.gate.n82 sg13g2_Clamp_N43N43D4R_0.gate.n80 0.853
R118 sg13g2_Clamp_N43N43D4R_0.gate.n110 sg13g2_Clamp_N43N43D4R_0.gate.n109 0.332192
R119 sg13g2_Clamp_N43N43D4R_0.gate.n111 sg13g2_Clamp_N43N43D4R_0.gate.n110 0.119159
R120 sg13g2_Clamp_N43N43D4R_0.gate sg13g2_Clamp_N43N43D4R_0.gate.n111 0.0570714
R121 sg13g2_Clamp_N43N43D4R_0.gate.n87 sg13g2_Clamp_N43N43D4R_0.gate.n86 0.0233437
R122 sg13g2_Clamp_N43N43D4R_0.gate.n88 sg13g2_Clamp_N43N43D4R_0.gate.n87 0.0233437
R123 sg13g2_Clamp_N43N43D4R_0.gate.n89 sg13g2_Clamp_N43N43D4R_0.gate.n88 0.0233437
R124 sg13g2_Clamp_N43N43D4R_0.gate.n90 sg13g2_Clamp_N43N43D4R_0.gate.n89 0.0233437
R125 sg13g2_Clamp_N43N43D4R_0.gate.n91 sg13g2_Clamp_N43N43D4R_0.gate.n90 0.0233437
R126 sg13g2_Clamp_N43N43D4R_0.gate.n92 sg13g2_Clamp_N43N43D4R_0.gate.n91 0.0233437
R127 sg13g2_Clamp_N43N43D4R_0.gate.n93 sg13g2_Clamp_N43N43D4R_0.gate.n92 0.0233437
R128 sg13g2_Clamp_N43N43D4R_0.gate.n94 sg13g2_Clamp_N43N43D4R_0.gate.n93 0.0233437
R129 sg13g2_Clamp_N43N43D4R_0.gate.n95 sg13g2_Clamp_N43N43D4R_0.gate.n94 0.0233437
R130 sg13g2_Clamp_N43N43D4R_0.gate.n96 sg13g2_Clamp_N43N43D4R_0.gate.n95 0.0233437
R131 sg13g2_Clamp_N43N43D4R_0.gate.n97 sg13g2_Clamp_N43N43D4R_0.gate.n96 0.0233437
R132 sg13g2_Clamp_N43N43D4R_0.gate.n98 sg13g2_Clamp_N43N43D4R_0.gate.n97 0.0233437
R133 sg13g2_Clamp_N43N43D4R_0.gate.n99 sg13g2_Clamp_N43N43D4R_0.gate.n98 0.0233437
R134 sg13g2_Clamp_N43N43D4R_0.gate.n100 sg13g2_Clamp_N43N43D4R_0.gate.n99 0.0233437
R135 sg13g2_Clamp_N43N43D4R_0.gate.n101 sg13g2_Clamp_N43N43D4R_0.gate.n100 0.0233437
R136 sg13g2_Clamp_N43N43D4R_0.gate.n102 sg13g2_Clamp_N43N43D4R_0.gate.n101 0.0233437
R137 sg13g2_Clamp_N43N43D4R_0.gate.n103 sg13g2_Clamp_N43N43D4R_0.gate.n102 0.0233437
R138 sg13g2_Clamp_N43N43D4R_0.gate.n104 sg13g2_Clamp_N43N43D4R_0.gate.n103 0.0233437
R139 sg13g2_Clamp_N43N43D4R_0.gate.n105 sg13g2_Clamp_N43N43D4R_0.gate.n104 0.0233437
R140 sg13g2_Clamp_N43N43D4R_0.gate.n106 sg13g2_Clamp_N43N43D4R_0.gate.n105 0.0233437
R141 sg13g2_Clamp_N43N43D4R_0.gate.n107 sg13g2_Clamp_N43N43D4R_0.gate.n106 0.0233437
R142 sg13g2_Clamp_N43N43D4R_0.gate.n108 sg13g2_Clamp_N43N43D4R_0.gate.n107 0.0233437
R143 sg13g2_Clamp_N43N43D4R_0.gate.n109 sg13g2_Clamp_N43N43D4R_0.gate.n108 0.0233437
R144 sg13g2_Clamp_N43N43D4R_0.gate.n83 sg13g2_Clamp_N43N43D4R_0.gate.t76 0.001
R145 sg13g2_Clamp_N43N43D4R_0.gate.n83 sg13g2_Clamp_N43N43D4R_0.gate.t114 0.001
R146 sg13g2_Clamp_N43N43D4R_0.gate.n0 sg13g2_Clamp_N43N43D4R_0.gate.t66 0.001
R147 sg13g2_Clamp_N43N43D4R_0.gate.n0 sg13g2_Clamp_N43N43D4R_0.gate.t109 0.001
R148 sg13g2_Clamp_N43N43D4R_0.gate.n1 sg13g2_Clamp_N43N43D4R_0.gate.t70 0.001
R149 sg13g2_Clamp_N43N43D4R_0.gate.n1 sg13g2_Clamp_N43N43D4R_0.gate.t85 0.001
R150 sg13g2_Clamp_N43N43D4R_0.gate.n3 sg13g2_Clamp_N43N43D4R_0.gate.t88 0.001
R151 sg13g2_Clamp_N43N43D4R_0.gate.n3 sg13g2_Clamp_N43N43D4R_0.gate.t32 0.001
R152 sg13g2_Clamp_N43N43D4R_0.gate.n5 sg13g2_Clamp_N43N43D4R_0.gate.t37 0.001
R153 sg13g2_Clamp_N43N43D4R_0.gate.n5 sg13g2_Clamp_N43N43D4R_0.gate.t99 0.001
R154 sg13g2_Clamp_N43N43D4R_0.gate.n7 sg13g2_Clamp_N43N43D4R_0.gate.t51 0.001
R155 sg13g2_Clamp_N43N43D4R_0.gate.n7 sg13g2_Clamp_N43N43D4R_0.gate.t68 0.001
R156 sg13g2_Clamp_N43N43D4R_0.gate.n9 sg13g2_Clamp_N43N43D4R_0.gate.t60 0.001
R157 sg13g2_Clamp_N43N43D4R_0.gate.n9 sg13g2_Clamp_N43N43D4R_0.gate.t103 0.001
R158 sg13g2_Clamp_N43N43D4R_0.gate.n11 sg13g2_Clamp_N43N43D4R_0.gate.t75 0.001
R159 sg13g2_Clamp_N43N43D4R_0.gate.n11 sg13g2_Clamp_N43N43D4R_0.gate.t89 0.001
R160 sg13g2_Clamp_N43N43D4R_0.gate.n13 sg13g2_Clamp_N43N43D4R_0.gate.t98 0.001
R161 sg13g2_Clamp_N43N43D4R_0.gate.n13 sg13g2_Clamp_N43N43D4R_0.gate.t47 0.001
R162 sg13g2_Clamp_N43N43D4R_0.gate.n15 sg13g2_Clamp_N43N43D4R_0.gate.t58 0.001
R163 sg13g2_Clamp_N43N43D4R_0.gate.n15 sg13g2_Clamp_N43N43D4R_0.gate.t72 0.001
R164 sg13g2_Clamp_N43N43D4R_0.gate.n17 sg13g2_Clamp_N43N43D4R_0.gate.t53 0.001
R165 sg13g2_Clamp_N43N43D4R_0.gate.n17 sg13g2_Clamp_N43N43D4R_0.gate.t69 0.001
R166 sg13g2_Clamp_N43N43D4R_0.gate.n19 sg13g2_Clamp_N43N43D4R_0.gate.t45 0.001
R167 sg13g2_Clamp_N43N43D4R_0.gate.n19 sg13g2_Clamp_N43N43D4R_0.gate.t106 0.001
R168 sg13g2_Clamp_N43N43D4R_0.gate.n21 sg13g2_Clamp_N43N43D4R_0.gate.t36 0.001
R169 sg13g2_Clamp_N43N43D4R_0.gate.n21 sg13g2_Clamp_N43N43D4R_0.gate.t50 0.001
R170 sg13g2_Clamp_N43N43D4R_0.gate.n23 sg13g2_Clamp_N43N43D4R_0.gate.t67 0.001
R171 sg13g2_Clamp_N43N43D4R_0.gate.n23 sg13g2_Clamp_N43N43D4R_0.gate.t110 0.001
R172 sg13g2_Clamp_N43N43D4R_0.gate.n25 sg13g2_Clamp_N43N43D4R_0.gate.t56 0.001
R173 sg13g2_Clamp_N43N43D4R_0.gate.n25 sg13g2_Clamp_N43N43D4R_0.gate.t102 0.001
R174 sg13g2_Clamp_N43N43D4R_0.gate.n27 sg13g2_Clamp_N43N43D4R_0.gate.t33 0.001
R175 sg13g2_Clamp_N43N43D4R_0.gate.n27 sg13g2_Clamp_N43N43D4R_0.gate.t49 0.001
R176 sg13g2_Clamp_N43N43D4R_0.gate.n29 sg13g2_Clamp_N43N43D4R_0.gate.t34 0.001
R177 sg13g2_Clamp_N43N43D4R_0.gate.n29 sg13g2_Clamp_N43N43D4R_0.gate.t105 0.001
R178 sg13g2_Clamp_N43N43D4R_0.gate.n31 sg13g2_Clamp_N43N43D4R_0.gate.t86 0.001
R179 sg13g2_Clamp_N43N43D4R_0.gate.n31 sg13g2_Clamp_N43N43D4R_0.gate.t96 0.001
R180 sg13g2_Clamp_N43N43D4R_0.gate.n33 sg13g2_Clamp_N43N43D4R_0.gate.t41 0.001
R181 sg13g2_Clamp_N43N43D4R_0.gate.n33 sg13g2_Clamp_N43N43D4R_0.gate.t55 0.001
R182 sg13g2_Clamp_N43N43D4R_0.gate.n35 sg13g2_Clamp_N43N43D4R_0.gate.t65 0.001
R183 sg13g2_Clamp_N43N43D4R_0.gate.n35 sg13g2_Clamp_N43N43D4R_0.gate.t82 0.001
R184 sg13g2_Clamp_N43N43D4R_0.gate.n37 sg13g2_Clamp_N43N43D4R_0.gate.t62 0.001
R185 sg13g2_Clamp_N43N43D4R_0.gate.n37 sg13g2_Clamp_N43N43D4R_0.gate.t78 0.001
R186 sg13g2_Clamp_N43N43D4R_0.gate.n39 sg13g2_Clamp_N43N43D4R_0.gate.t54 0.001
R187 sg13g2_Clamp_N43N43D4R_0.gate.n39 sg13g2_Clamp_N43N43D4R_0.gate.t108 0.001
R188 sg13g2_Clamp_N43N43D4R_0.gate.n41 sg13g2_Clamp_N43N43D4R_0.gate.t46 0.001
R189 sg13g2_Clamp_N43N43D4R_0.gate.n41 sg13g2_Clamp_N43N43D4R_0.gate.t61 0.001
R190 sg13g2_Clamp_N43N43D4R_0.gate.n43 sg13g2_Clamp_N43N43D4R_0.gate.t77 0.001
R191 sg13g2_Clamp_N43N43D4R_0.gate.n43 sg13g2_Clamp_N43N43D4R_0.gate.t115 0.001
R192 sg13g2_Clamp_N43N43D4R_0.gate.n45 sg13g2_Clamp_N43N43D4R_0.gate.t31 0.001
R193 sg13g2_Clamp_N43N43D4R_0.gate.n45 sg13g2_Clamp_N43N43D4R_0.gate.t104 0.001
R194 sg13g2_Clamp_N43N43D4R_0.gate.n47 sg13g2_Clamp_N43N43D4R_0.gate.t42 0.001
R195 sg13g2_Clamp_N43N43D4R_0.gate.n47 sg13g2_Clamp_N43N43D4R_0.gate.t57 0.001
R196 sg13g2_Clamp_N43N43D4R_0.gate.n49 sg13g2_Clamp_N43N43D4R_0.gate.t48 0.001
R197 sg13g2_Clamp_N43N43D4R_0.gate.n49 sg13g2_Clamp_N43N43D4R_0.gate.t101 0.001
R198 sg13g2_Clamp_N43N43D4R_0.gate.n51 sg13g2_Clamp_N43N43D4R_0.gate.t63 0.001
R199 sg13g2_Clamp_N43N43D4R_0.gate.n51 sg13g2_Clamp_N43N43D4R_0.gate.t80 0.001
R200 sg13g2_Clamp_N43N43D4R_0.gate.n53 sg13g2_Clamp_N43N43D4R_0.gate.t90 0.001
R201 sg13g2_Clamp_N43N43D4R_0.gate.n53 sg13g2_Clamp_N43N43D4R_0.gate.t35 0.001
R202 sg13g2_Clamp_N43N43D4R_0.gate.n55 sg13g2_Clamp_N43N43D4R_0.gate.t87 0.001
R203 sg13g2_Clamp_N43N43D4R_0.gate.n55 sg13g2_Clamp_N43N43D4R_0.gate.t97 0.001
R204 sg13g2_Clamp_N43N43D4R_0.gate.n57 sg13g2_Clamp_N43N43D4R_0.gate.t43 0.001
R205 sg13g2_Clamp_N43N43D4R_0.gate.n57 sg13g2_Clamp_N43N43D4R_0.gate.t59 0.001
R206 sg13g2_Clamp_N43N43D4R_0.gate.n59 sg13g2_Clamp_N43N43D4R_0.gate.t74 0.001
R207 sg13g2_Clamp_N43N43D4R_0.gate.n59 sg13g2_Clamp_N43N43D4R_0.gate.t112 0.001
R208 sg13g2_Clamp_N43N43D4R_0.gate.n61 sg13g2_Clamp_N43N43D4R_0.gate.t92 0.001
R209 sg13g2_Clamp_N43N43D4R_0.gate.n61 sg13g2_Clamp_N43N43D4R_0.gate.t39 0.001
R210 sg13g2_Clamp_N43N43D4R_0.gate.n63 sg13g2_Clamp_N43N43D4R_0.gate.t93 0.001
R211 sg13g2_Clamp_N43N43D4R_0.gate.n63 sg13g2_Clamp_N43N43D4R_0.gate.t40 0.001
R212 sg13g2_Clamp_N43N43D4R_0.gate.n65 sg13g2_Clamp_N43N43D4R_0.gate.t44 0.001
R213 sg13g2_Clamp_N43N43D4R_0.gate.n65 sg13g2_Clamp_N43N43D4R_0.gate.t100 0.001
R214 sg13g2_Clamp_N43N43D4R_0.gate.n67 sg13g2_Clamp_N43N43D4R_0.gate.t79 0.001
R215 sg13g2_Clamp_N43N43D4R_0.gate.n67 sg13g2_Clamp_N43N43D4R_0.gate.t116 0.001
R216 sg13g2_Clamp_N43N43D4R_0.gate.n69 sg13g2_Clamp_N43N43D4R_0.gate.t83 0.001
R217 sg13g2_Clamp_N43N43D4R_0.gate.n69 sg13g2_Clamp_N43N43D4R_0.gate.t94 0.001
R218 sg13g2_Clamp_N43N43D4R_0.gate.n71 sg13g2_Clamp_N43N43D4R_0.gate.t84 0.001
R219 sg13g2_Clamp_N43N43D4R_0.gate.n71 sg13g2_Clamp_N43N43D4R_0.gate.t95 0.001
R220 sg13g2_Clamp_N43N43D4R_0.gate.n73 sg13g2_Clamp_N43N43D4R_0.gate.t71 0.001
R221 sg13g2_Clamp_N43N43D4R_0.gate.n73 sg13g2_Clamp_N43N43D4R_0.gate.t111 0.001
R222 sg13g2_Clamp_N43N43D4R_0.gate.n75 sg13g2_Clamp_N43N43D4R_0.gate.t64 0.001
R223 sg13g2_Clamp_N43N43D4R_0.gate.n75 sg13g2_Clamp_N43N43D4R_0.gate.t81 0.001
R224 sg13g2_Clamp_N43N43D4R_0.gate.n77 sg13g2_Clamp_N43N43D4R_0.gate.t91 0.001
R225 sg13g2_Clamp_N43N43D4R_0.gate.n77 sg13g2_Clamp_N43N43D4R_0.gate.t38 0.001
R226 sg13g2_Clamp_N43N43D4R_0.gate.n79 sg13g2_Clamp_N43N43D4R_0.gate.t52 0.001
R227 sg13g2_Clamp_N43N43D4R_0.gate.n79 sg13g2_Clamp_N43N43D4R_0.gate.t107 0.001
R228 sg13g2_Clamp_N43N43D4R_0.gate.n81 sg13g2_Clamp_N43N43D4R_0.gate.t73 0.001
R229 sg13g2_Clamp_N43N43D4R_0.gate.n81 sg13g2_Clamp_N43N43D4R_0.gate.t113 0.001
R230 iovdd.n625 iovdd.n109 25.498
R231 iovdd.n604 iovdd.n603 9.7146
R232 iovdd.n400 iovdd.n399 9.7146
R233 iovdd.n391 iovdd.n390 9.7146
R234 iovdd.n377 iovdd.n376 9.7146
R235 iovdd.n367 iovdd.n366 9.7146
R236 iovdd.n353 iovdd.n352 9.7146
R237 iovdd.n343 iovdd.n342 9.7146
R238 iovdd.n330 iovdd.n329 9.7146
R239 iovdd.n313 iovdd.n312 9.7146
R240 iovdd.n305 iovdd.n304 9.7146
R241 iovdd.n296 iovdd.n295 9.7146
R242 iovdd.n282 iovdd.n281 9.7146
R243 iovdd.n272 iovdd.n271 9.7146
R244 iovdd.n258 iovdd.n257 9.7146
R245 iovdd.n248 iovdd.n247 9.7146
R246 iovdd.n235 iovdd.n234 9.7146
R247 iovdd.n220 iovdd.n219 9.7146
R248 iovdd.n211 iovdd.n210 9.7146
R249 iovdd.n204 iovdd.n203 9.7146
R250 iovdd.n159 iovdd.n158 9.7146
R251 iovdd.n168 iovdd.n167 9.7146
R252 iovdd.n609 iovdd.n608 9.7146
R253 iovdd.n109 iovdd.t88 4.97569
R254 iovdd.n143 iovdd.n140 4.5146
R255 iovdd.n627 iovdd.n626 4.5005
R256 iovdd.n111 iovdd.n107 4.5005
R257 iovdd.n409 iovdd.n408 4.5005
R258 iovdd.n407 iovdd.n405 4.5005
R259 iovdd.n406 iovdd.n396 4.5005
R260 iovdd.n433 iovdd.n373 4.5005
R261 iovdd.n441 iovdd.n440 4.5005
R262 iovdd.n443 iovdd.n442 4.5005
R263 iovdd.n451 iovdd.n349 4.5005
R264 iovdd.n459 iovdd.n458 4.5005
R265 iovdd.n461 iovdd.n460 4.5005
R266 iovdd.n469 iovdd.n326 4.5005
R267 iovdd.n477 iovdd.n476 4.5005
R268 iovdd.n479 iovdd.n478 4.5005
R269 iovdd.n324 iovdd.n318 4.5005
R270 iovdd.n323 iovdd.n310 4.5005
R271 iovdd.n322 iovdd.n301 4.5005
R272 iovdd.n508 iovdd.n278 4.5005
R273 iovdd.n516 iovdd.n515 4.5005
R274 iovdd.n518 iovdd.n517 4.5005
R275 iovdd.n526 iovdd.n254 4.5005
R276 iovdd.n534 iovdd.n533 4.5005
R277 iovdd.n536 iovdd.n535 4.5005
R278 iovdd.n544 iovdd.n231 4.5005
R279 iovdd.n552 iovdd.n551 4.5005
R280 iovdd.n555 iovdd.n554 4.5005
R281 iovdd.n230 iovdd.n225 4.5005
R282 iovdd.n229 iovdd.n216 4.5005
R283 iovdd.n576 iovdd.n153 4.5005
R284 iovdd.n585 iovdd.n584 4.5005
R285 iovdd.n192 iovdd.n152 4.5005
R286 iovdd.n185 iovdd.n184 4.5005
R287 iovdd.n176 iovdd.n144 4.5005
R288 iovdd.n596 iovdd.n595 4.5005
R289 iovdd.n145 iovdd.n143 4.5005
R290 iovdd.n595 iovdd.n594 4.5005
R291 iovdd.n146 iovdd.n144 4.5005
R292 iovdd.n184 iovdd.n151 4.5005
R293 iovdd.n587 iovdd.n152 4.5005
R294 iovdd.n586 iovdd.n585 4.5005
R295 iovdd.n153 iovdd.n78 4.5005
R296 iovdd.n229 iovdd.n79 4.5005
R297 iovdd.n230 iovdd.n80 4.5005
R298 iovdd.n554 iovdd.n553 4.5005
R299 iovdd.n552 iovdd.n83 4.5005
R300 iovdd.n231 iovdd.n84 4.5005
R301 iovdd.n535 iovdd.n85 4.5005
R302 iovdd.n534 iovdd.n86 4.5005
R303 iovdd.n254 iovdd.n87 4.5005
R304 iovdd.n517 iovdd.n88 4.5005
R305 iovdd.n516 iovdd.n89 4.5005
R306 iovdd.n278 iovdd.n90 4.5005
R307 iovdd.n322 iovdd.n91 4.5005
R308 iovdd.n323 iovdd.n92 4.5005
R309 iovdd.n324 iovdd.n93 4.5005
R310 iovdd.n478 iovdd.n94 4.5005
R311 iovdd.n477 iovdd.n95 4.5005
R312 iovdd.n326 iovdd.n325 4.5005
R313 iovdd.n460 iovdd.n97 4.5005
R314 iovdd.n459 iovdd.n98 4.5005
R315 iovdd.n349 iovdd.n99 4.5005
R316 iovdd.n442 iovdd.n100 4.5005
R317 iovdd.n441 iovdd.n101 4.5005
R318 iovdd.n373 iovdd.n102 4.5005
R319 iovdd.n406 iovdd.n103 4.5005
R320 iovdd.n407 iovdd.n104 4.5005
R321 iovdd.n408 iovdd.n105 4.5005
R322 iovdd.n107 iovdd.n106 4.5005
R323 iovdd.n628 iovdd.n627 4.5005
R324 iovdd.n804 iovdd.n754 3.31474
R325 iovdd.n804 iovdd.n758 3.31474
R326 iovdd.n804 iovdd.n764 3.31474
R327 iovdd.n804 iovdd.n768 3.31474
R328 iovdd.n804 iovdd.n774 3.31474
R329 iovdd.n804 iovdd.n778 3.31474
R330 iovdd.n804 iovdd.n782 3.31474
R331 iovdd.n804 iovdd.n788 3.31474
R332 iovdd.n804 iovdd.n792 3.31474
R333 iovdd.n804 iovdd.n798 3.31474
R334 iovdd.n804 iovdd.n803 3.31474
R335 iovdd.n804 iovdd.n756 3.31457
R336 iovdd.n804 iovdd.n760 3.31457
R337 iovdd.n804 iovdd.n766 3.31457
R338 iovdd.n804 iovdd.n770 3.31457
R339 iovdd.n804 iovdd.n776 3.31457
R340 iovdd.n804 iovdd.n780 3.31457
R341 iovdd.n804 iovdd.n786 3.31457
R342 iovdd.n804 iovdd.n790 3.31457
R343 iovdd.n804 iovdd.n794 3.31457
R344 iovdd.n804 iovdd.n800 3.31457
R345 iovdd.n795 iovdd.t115 3.28171
R346 iovdd.n761 iovdd.t106 3.28171
R347 iovdd.n801 iovdd.t93 3.28171
R348 iovdd.n802 iovdd.t117 3.28171
R349 iovdd.n799 iovdd.t109 3.28171
R350 iovdd.n797 iovdd.t122 3.28171
R351 iovdd.n793 iovdd.t113 3.28171
R352 iovdd.n791 iovdd.t95 3.28171
R353 iovdd.n789 iovdd.t101 3.28171
R354 iovdd.n787 iovdd.t94 3.28171
R355 iovdd.n785 iovdd.t108 3.28171
R356 iovdd.n783 iovdd.t98 3.28171
R357 iovdd.n781 iovdd.t111 3.28171
R358 iovdd.n779 iovdd.t92 3.28171
R359 iovdd.n777 iovdd.t103 3.28171
R360 iovdd.n775 iovdd.t96 3.28171
R361 iovdd.n773 iovdd.t105 3.28171
R362 iovdd.n771 iovdd.t99 3.28171
R363 iovdd.n769 iovdd.t100 3.28171
R364 iovdd.n767 iovdd.t90 3.28171
R365 iovdd.n765 iovdd.t104 3.28171
R366 iovdd.n763 iovdd.t97 3.28171
R367 iovdd.n759 iovdd.t131 3.28171
R368 iovdd.n757 iovdd.t102 3.28171
R369 iovdd.n755 iovdd.t91 3.28171
R370 iovdd.n753 iovdd.t114 3.28171
R371 iovdd.n804 iovdd.n784 2.73027
R372 iovdd.n804 iovdd.n762 2.73011
R373 iovdd.n804 iovdd.n772 2.73011
R374 iovdd.n804 iovdd.n796 2.73011
R375 iovdd.n630 iovdd.n628 2.2005
R376 iovdd.n631 iovdd.n106 2.2005
R377 iovdd.n632 iovdd.n105 2.2005
R378 iovdd.n634 iovdd.n104 2.2005
R379 iovdd.n635 iovdd.n103 2.2005
R380 iovdd.n637 iovdd.n102 2.2005
R381 iovdd.n638 iovdd.n101 2.2005
R382 iovdd.n640 iovdd.n100 2.2005
R383 iovdd.n641 iovdd.n99 2.2005
R384 iovdd.n643 iovdd.n98 2.2005
R385 iovdd.n644 iovdd.n97 2.2005
R386 iovdd.n325 iovdd.n96 2.2005
R387 iovdd.n648 iovdd.n95 2.2005
R388 iovdd.n649 iovdd.n94 2.2005
R389 iovdd.n651 iovdd.n93 2.2005
R390 iovdd.n652 iovdd.n92 2.2005
R391 iovdd.n654 iovdd.n91 2.2005
R392 iovdd.n655 iovdd.n90 2.2005
R393 iovdd.n657 iovdd.n89 2.2005
R394 iovdd.n658 iovdd.n88 2.2005
R395 iovdd.n660 iovdd.n87 2.2005
R396 iovdd.n661 iovdd.n86 2.2005
R397 iovdd.n663 iovdd.n85 2.2005
R398 iovdd.n664 iovdd.n84 2.2005
R399 iovdd.n665 iovdd.n83 2.2005
R400 iovdd.n553 iovdd.n81 2.2005
R401 iovdd.n670 iovdd.n80 2.2005
R402 iovdd.n671 iovdd.n79 2.2005
R403 iovdd.n672 iovdd.n78 2.2005
R404 iovdd.n586 iovdd.n77 2.2005
R405 iovdd.n588 iovdd.n587 2.2005
R406 iovdd.n589 iovdd.n151 2.2005
R407 iovdd.n148 iovdd.n146 2.2005
R408 iovdd.n594 iovdd.n593 2.2005
R409 iovdd.n147 iovdd.n145 2.2005
R410 iovdd.n400 iovdd.t59 1.78531
R411 iovdd.n401 iovdd.t78 1.78531
R412 iovdd.n402 iovdd.t7 1.78531
R413 iovdd.n403 iovdd.t33 1.78531
R414 iovdd.n391 iovdd.t21 1.78531
R415 iovdd.n392 iovdd.t51 1.78531
R416 iovdd.n393 iovdd.t31 1.78531
R417 iovdd.n394 iovdd.t15 1.78531
R418 iovdd.n377 iovdd.t3 1.78531
R419 iovdd.n378 iovdd.t40 1.78531
R420 iovdd.n379 iovdd.t81 1.78531
R421 iovdd.n380 iovdd.t75 1.78531
R422 iovdd.n367 iovdd.t69 1.78531
R423 iovdd.n368 iovdd.t18 1.78531
R424 iovdd.n369 iovdd.t24 1.78531
R425 iovdd.n370 iovdd.t8 1.78531
R426 iovdd.n353 iovdd.t55 1.78531
R427 iovdd.n354 iovdd.t77 1.78531
R428 iovdd.n355 iovdd.t4 1.78531
R429 iovdd.n356 iovdd.t87 1.78531
R430 iovdd.n343 iovdd.t43 1.78531
R431 iovdd.n344 iovdd.t67 1.78531
R432 iovdd.n345 iovdd.t29 1.78531
R433 iovdd.n346 iovdd.t14 1.78531
R434 iovdd.n330 iovdd.t2 1.78531
R435 iovdd.n331 iovdd.t34 1.78531
R436 iovdd.n332 iovdd.t10 1.78531
R437 iovdd.n333 iovdd.t74 1.78531
R438 iovdd.n313 iovdd.t23 1.78531
R439 iovdd.n314 iovdd.t16 1.78531
R440 iovdd.n315 iovdd.t73 1.78531
R441 iovdd.n316 iovdd.t63 1.78531
R442 iovdd.n305 iovdd.t44 1.78531
R443 iovdd.n306 iovdd.t66 1.78531
R444 iovdd.n307 iovdd.t62 1.78531
R445 iovdd.n308 iovdd.t50 1.78531
R446 iovdd.n296 iovdd.t42 1.78531
R447 iovdd.n297 iovdd.t64 1.78531
R448 iovdd.n298 iovdd.t26 1.78531
R449 iovdd.n299 iovdd.t9 1.78531
R450 iovdd.n282 iovdd.t25 1.78531
R451 iovdd.n283 iovdd.t53 1.78531
R452 iovdd.n284 iovdd.t45 1.78531
R453 iovdd.n285 iovdd.t32 1.78531
R454 iovdd.n272 iovdd.t20 1.78531
R455 iovdd.n273 iovdd.t49 1.78531
R456 iovdd.n274 iovdd.t86 1.78531
R457 iovdd.n275 iovdd.t82 1.78531
R458 iovdd.n258 iovdd.t1 1.78531
R459 iovdd.n259 iovdd.t38 1.78531
R460 iovdd.n260 iovdd.t61 1.78531
R461 iovdd.n261 iovdd.t47 1.78531
R462 iovdd.n248 iovdd.t52 1.78531
R463 iovdd.n249 iovdd.t6 1.78531
R464 iovdd.n250 iovdd.t68 1.78531
R465 iovdd.n251 iovdd.t58 1.78531
R466 iovdd.n235 iovdd.t48 1.78531
R467 iovdd.n236 iovdd.t72 1.78531
R468 iovdd.n237 iovdd.t37 1.78531
R469 iovdd.n238 iovdd.t19 1.78531
R470 iovdd.n220 iovdd.t36 1.78531
R471 iovdd.n221 iovdd.t60 1.78531
R472 iovdd.n222 iovdd.t54 1.78531
R473 iovdd.n223 iovdd.t41 1.78531
R474 iovdd.n211 iovdd.t30 1.78531
R475 iovdd.n212 iovdd.t56 1.78531
R476 iovdd.n213 iovdd.t0 1.78531
R477 iovdd.n214 iovdd.t84 1.78531
R478 iovdd.n204 iovdd.t12 1.78531
R479 iovdd.n205 iovdd.t5 1.78531
R480 iovdd.n206 iovdd.t65 1.78531
R481 iovdd.n207 iovdd.t57 1.78531
R482 iovdd.n159 iovdd.t35 1.78531
R483 iovdd.n160 iovdd.t28 1.78531
R484 iovdd.n161 iovdd.t79 1.78531
R485 iovdd.n162 iovdd.t71 1.78531
R486 iovdd.n168 iovdd.t17 1.78531
R487 iovdd.n169 iovdd.t46 1.78531
R488 iovdd.n170 iovdd.t13 1.78531
R489 iovdd.n171 iovdd.t80 1.78531
R490 iovdd.n609 iovdd.t70 1.78531
R491 iovdd.n610 iovdd.t83 1.78531
R492 iovdd.n611 iovdd.t27 1.78531
R493 iovdd.n612 iovdd.t11 1.78531
R494 iovdd.n603 iovdd.t76 1.78502
R495 iovdd.n602 iovdd.t85 1.78502
R496 iovdd.n601 iovdd.t39 1.78502
R497 iovdd.n600 iovdd.t22 1.78502
R498 iovdd.n624 iovdd.n108 1.5005
R499 iovdd.n623 iovdd.n622 1.5005
R500 iovdd.n621 iovdd.n110 1.5005
R501 iovdd.n620 iovdd.n619 1.5005
R502 iovdd.n618 iovdd.n617 1.5005
R503 iovdd.n616 iovdd.n112 1.5005
R504 iovdd.n615 iovdd.n614 1.5005
R505 iovdd.n114 iovdd.n113 1.5005
R506 iovdd.n411 iovdd.n410 1.5005
R507 iovdd.n413 iovdd.n412 1.5005
R508 iovdd.n414 iovdd.n404 1.5005
R509 iovdd.n416 iovdd.n415 1.5005
R510 iovdd.n418 iovdd.n398 1.5005
R511 iovdd.n420 iovdd.n419 1.5005
R512 iovdd.n421 iovdd.n397 1.5005
R513 iovdd.n423 iovdd.n422 1.5005
R514 iovdd.n425 iovdd.n424 1.5005
R515 iovdd.n426 iovdd.n395 1.5005
R516 iovdd.n428 iovdd.n427 1.5005
R517 iovdd.n430 iovdd.n389 1.5005
R518 iovdd.n432 iovdd.n431 1.5005
R519 iovdd.n434 iovdd.n388 1.5005
R520 iovdd.n436 iovdd.n435 1.5005
R521 iovdd.n437 iovdd.n375 1.5005
R522 iovdd.n439 iovdd.n438 1.5005
R523 iovdd.n386 iovdd.n374 1.5005
R524 iovdd.n385 iovdd.n384 1.5005
R525 iovdd.n383 iovdd.n382 1.5005
R526 iovdd.n381 iovdd.n372 1.5005
R527 iovdd.n444 iovdd.n371 1.5005
R528 iovdd.n446 iovdd.n445 1.5005
R529 iovdd.n448 iovdd.n365 1.5005
R530 iovdd.n450 iovdd.n449 1.5005
R531 iovdd.n452 iovdd.n364 1.5005
R532 iovdd.n454 iovdd.n453 1.5005
R533 iovdd.n455 iovdd.n351 1.5005
R534 iovdd.n457 iovdd.n456 1.5005
R535 iovdd.n362 iovdd.n350 1.5005
R536 iovdd.n361 iovdd.n360 1.5005
R537 iovdd.n359 iovdd.n358 1.5005
R538 iovdd.n357 iovdd.n348 1.5005
R539 iovdd.n462 iovdd.n347 1.5005
R540 iovdd.n464 iovdd.n463 1.5005
R541 iovdd.n466 iovdd.n341 1.5005
R542 iovdd.n468 iovdd.n467 1.5005
R543 iovdd.n470 iovdd.n340 1.5005
R544 iovdd.n472 iovdd.n471 1.5005
R545 iovdd.n473 iovdd.n328 1.5005
R546 iovdd.n475 iovdd.n474 1.5005
R547 iovdd.n338 iovdd.n327 1.5005
R548 iovdd.n337 iovdd.n336 1.5005
R549 iovdd.n335 iovdd.n334 1.5005
R550 iovdd.n321 iovdd.n320 1.5005
R551 iovdd.n481 iovdd.n480 1.5005
R552 iovdd.n482 iovdd.n319 1.5005
R553 iovdd.n484 iovdd.n483 1.5005
R554 iovdd.n486 iovdd.n485 1.5005
R555 iovdd.n487 iovdd.n311 1.5005
R556 iovdd.n489 iovdd.n488 1.5005
R557 iovdd.n490 iovdd.n309 1.5005
R558 iovdd.n492 iovdd.n491 1.5005
R559 iovdd.n493 iovdd.n303 1.5005
R560 iovdd.n496 iovdd.n495 1.5005
R561 iovdd.n497 iovdd.n302 1.5005
R562 iovdd.n499 iovdd.n498 1.5005
R563 iovdd.n501 iovdd.n500 1.5005
R564 iovdd.n502 iovdd.n300 1.5005
R565 iovdd.n504 iovdd.n503 1.5005
R566 iovdd.n506 iovdd.n294 1.5005
R567 iovdd.n508 iovdd.n507 1.5005
R568 iovdd.n509 iovdd.n293 1.5005
R569 iovdd.n511 iovdd.n510 1.5005
R570 iovdd.n512 iovdd.n280 1.5005
R571 iovdd.n514 iovdd.n513 1.5005
R572 iovdd.n291 iovdd.n279 1.5005
R573 iovdd.n290 iovdd.n289 1.5005
R574 iovdd.n288 iovdd.n287 1.5005
R575 iovdd.n286 iovdd.n277 1.5005
R576 iovdd.n519 iovdd.n276 1.5005
R577 iovdd.n521 iovdd.n520 1.5005
R578 iovdd.n523 iovdd.n270 1.5005
R579 iovdd.n525 iovdd.n524 1.5005
R580 iovdd.n527 iovdd.n269 1.5005
R581 iovdd.n529 iovdd.n528 1.5005
R582 iovdd.n530 iovdd.n256 1.5005
R583 iovdd.n532 iovdd.n531 1.5005
R584 iovdd.n267 iovdd.n255 1.5005
R585 iovdd.n266 iovdd.n265 1.5005
R586 iovdd.n264 iovdd.n263 1.5005
R587 iovdd.n262 iovdd.n253 1.5005
R588 iovdd.n537 iovdd.n252 1.5005
R589 iovdd.n539 iovdd.n538 1.5005
R590 iovdd.n540 iovdd.n246 1.5005
R591 iovdd.n543 iovdd.n542 1.5005
R592 iovdd.n545 iovdd.n245 1.5005
R593 iovdd.n547 iovdd.n546 1.5005
R594 iovdd.n548 iovdd.n233 1.5005
R595 iovdd.n550 iovdd.n549 1.5005
R596 iovdd.n244 iovdd.n232 1.5005
R597 iovdd.n242 iovdd.n241 1.5005
R598 iovdd.n240 iovdd.n239 1.5005
R599 iovdd.n228 iovdd.n227 1.5005
R600 iovdd.n557 iovdd.n556 1.5005
R601 iovdd.n558 iovdd.n226 1.5005
R602 iovdd.n560 iovdd.n559 1.5005
R603 iovdd.n562 iovdd.n561 1.5005
R604 iovdd.n563 iovdd.n218 1.5005
R605 iovdd.n565 iovdd.n564 1.5005
R606 iovdd.n566 iovdd.n217 1.5005
R607 iovdd.n568 iovdd.n567 1.5005
R608 iovdd.n570 iovdd.n569 1.5005
R609 iovdd.n572 iovdd.n571 1.5005
R610 iovdd.n573 iovdd.n209 1.5005
R611 iovdd.n575 iovdd.n574 1.5005
R612 iovdd.n577 iovdd.n208 1.5005
R613 iovdd.n579 iovdd.n578 1.5005
R614 iovdd.n580 iovdd.n155 1.5005
R615 iovdd.n583 iovdd.n582 1.5005
R616 iovdd.n202 iovdd.n154 1.5005
R617 iovdd.n201 iovdd.n200 1.5005
R618 iovdd.n199 iovdd.n156 1.5005
R619 iovdd.n198 iovdd.n197 1.5005
R620 iovdd.n196 iovdd.n157 1.5005
R621 iovdd.n194 iovdd.n193 1.5005
R622 iovdd.n191 iovdd.n163 1.5005
R623 iovdd.n190 iovdd.n189 1.5005
R624 iovdd.n188 iovdd.n164 1.5005
R625 iovdd.n187 iovdd.n186 1.5005
R626 iovdd.n183 iovdd.n165 1.5005
R627 iovdd.n182 iovdd.n181 1.5005
R628 iovdd.n179 iovdd.n166 1.5005
R629 iovdd.n178 iovdd.n177 1.5005
R630 iovdd.n175 iovdd.n172 1.5005
R631 iovdd.n174 iovdd.n173 1.5005
R632 iovdd.n142 iovdd.n141 1.5005
R633 iovdd.n598 iovdd.n597 1.5005
R634 iovdd.n138 iovdd.n116 1.49387
R635 iovdd.n139 iovdd.n138 1.45493
R636 iovdd.n139 iovdd.n137 1.45278
R637 iovdd.n137 iovdd.n116 1.41784
R638 iovdd.n806 iovdd.n805 1.41716
R639 iovdd.n806 iovdd.n750 1.37269
R640 iovdd.n805 iovdd.n751 1.35023
R641 iovdd.n801 iovdd.n750 1.34472
R642 iovdd.n752 iovdd.n751 1.2534
R643 iovdd.n753 iovdd.n752 1.19837
R644 iovdd.n149 iovdd.n147 1.106
R645 iovdd.n593 iovdd.n592 1.1005
R646 iovdd.n591 iovdd.n148 1.1005
R647 iovdd.n590 iovdd.n589 1.1005
R648 iovdd.n588 iovdd.n150 1.1005
R649 iovdd.n77 iovdd.n75 1.1005
R650 iovdd.n673 iovdd.n672 1.1005
R651 iovdd.n671 iovdd.n76 1.1005
R652 iovdd.n670 iovdd.n669 1.1005
R653 iovdd.n668 iovdd.n81 1.1005
R654 iovdd.n666 iovdd.n665 1.1005
R655 iovdd.n664 iovdd.n82 1.1005
R656 iovdd.n663 iovdd.n662 1.1005
R657 iovdd.n661 iovdd.n46 1.1005
R658 iovdd.n648 iovdd.n647 1.1005
R659 iovdd.n646 iovdd.n96 1.1005
R660 iovdd.n645 iovdd.n644 1.1005
R661 iovdd.n630 iovdd.n629 1.1005
R662 iovdd.n631 iovdd.n18 1.1005
R663 iovdd.n606 iovdd.n129 0.99443
R664 iovdd.n606 iovdd.n121 0.994252
R665 iovdd.n606 iovdd.n136 0.868409
R666 iovdd.n606 iovdd.n134 0.868409
R667 iovdd.n606 iovdd.n132 0.868409
R668 iovdd.n606 iovdd.n130 0.868409
R669 iovdd.n606 iovdd.n127 0.868409
R670 iovdd.n606 iovdd.n125 0.868409
R671 iovdd.n606 iovdd.n123 0.868409
R672 iovdd.n606 iovdd.n120 0.868409
R673 iovdd.n606 iovdd.n118 0.868409
R674 iovdd.n606 iovdd.n115 0.868254
R675 iovdd.n606 iovdd.n135 0.868254
R676 iovdd.n606 iovdd.n133 0.868254
R677 iovdd.n606 iovdd.n131 0.868254
R678 iovdd.n606 iovdd.n128 0.868254
R679 iovdd.n606 iovdd.n126 0.868254
R680 iovdd.n606 iovdd.n124 0.868254
R681 iovdd.n606 iovdd.n122 0.868254
R682 iovdd.n606 iovdd.n119 0.868254
R683 iovdd.n606 iovdd.n117 0.868254
R684 iovdd iovdd.n599 0.83073
R685 iovdd.n417 iovdd 0.83073
R686 iovdd.n429 iovdd 0.83073
R687 iovdd.n387 iovdd 0.83073
R688 iovdd.n447 iovdd 0.83073
R689 iovdd.n363 iovdd 0.83073
R690 iovdd.n465 iovdd 0.83073
R691 iovdd.n339 iovdd 0.83073
R692 iovdd.n317 iovdd 0.83073
R693 iovdd.n494 iovdd 0.83073
R694 iovdd.n505 iovdd 0.83073
R695 iovdd.n292 iovdd 0.83073
R696 iovdd.n522 iovdd 0.83073
R697 iovdd.n268 iovdd 0.83073
R698 iovdd.n541 iovdd 0.83073
R699 iovdd.n243 iovdd 0.83073
R700 iovdd.n224 iovdd 0.83073
R701 iovdd.n215 iovdd 0.83073
R702 iovdd.n581 iovdd 0.83073
R703 iovdd.n195 iovdd 0.83073
R704 iovdd.n180 iovdd 0.83073
R705 iovdd.n613 iovdd 0.83073
R706 iovdd.n693 iovdd.n690 0.826084
R707 iovdd.n1109 iovdd.n1108 0.826084
R708 iovdd.n970 iovdd.n966 0.826084
R709 iovdd.n867 iovdd.n866 0.822133
R710 iovdd.n866 iovdd.n865 0.818682
R711 iovdd.n864 iovdd.n862 0.818682
R712 iovdd.n874 iovdd.n861 0.818682
R713 iovdd.n875 iovdd.n860 0.818682
R714 iovdd.n859 iovdd.n857 0.818682
R715 iovdd.n858 iovdd.n848 0.818682
R716 iovdd.n885 iovdd.n847 0.818682
R717 iovdd.n886 iovdd.n846 0.818682
R718 iovdd.n845 iovdd.n843 0.818682
R719 iovdd.n844 iovdd.n836 0.818682
R720 iovdd.n896 iovdd.n835 0.818682
R721 iovdd.n897 iovdd.n834 0.818682
R722 iovdd.n833 iovdd.n831 0.818682
R723 iovdd.n832 iovdd.n823 0.818682
R724 iovdd.n907 iovdd.n822 0.818682
R725 iovdd.n908 iovdd.n821 0.818682
R726 iovdd.n820 iovdd.n818 0.818682
R727 iovdd.n819 iovdd.n809 0.818682
R728 iovdd.n918 iovdd.n808 0.818682
R729 iovdd.n919 iovdd.n807 0.818682
R730 iovdd.n749 iovdd.n745 0.818682
R731 iovdd.n928 iovdd.n744 0.818682
R732 iovdd.n929 iovdd.n743 0.818682
R733 iovdd.n742 iovdd.n740 0.818682
R734 iovdd.n741 iovdd.n732 0.818682
R735 iovdd.n939 iovdd.n731 0.818682
R736 iovdd.n940 iovdd.n730 0.818682
R737 iovdd.n729 iovdd.n727 0.818682
R738 iovdd.n728 iovdd.n719 0.818682
R739 iovdd.n950 iovdd.n718 0.818682
R740 iovdd.n951 iovdd.n717 0.818682
R741 iovdd.n716 iovdd.n680 0.818682
R742 iovdd.n715 iovdd.n714 0.818682
R743 iovdd.n682 iovdd.n681 0.818682
R744 iovdd.n703 iovdd.n702 0.818682
R745 iovdd.n701 iovdd.n689 0.818682
R746 iovdd.n700 iovdd.n699 0.818682
R747 iovdd.n692 iovdd.n691 0.818682
R748 iovdd.n699 iovdd.n698 0.818682
R749 iovdd.n689 iovdd.n687 0.818682
R750 iovdd.n704 iovdd.n703 0.818682
R751 iovdd.n683 iovdd.n682 0.818682
R752 iovdd.n714 iovdd.n713 0.818682
R753 iovdd.n680 iovdd.n678 0.818682
R754 iovdd.n952 iovdd.n951 0.818682
R755 iovdd.n950 iovdd.n949 0.818682
R756 iovdd.n720 iovdd.n719 0.818682
R757 iovdd.n727 iovdd.n725 0.818682
R758 iovdd.n941 iovdd.n940 0.818682
R759 iovdd.n939 iovdd.n938 0.818682
R760 iovdd.n733 iovdd.n732 0.818682
R761 iovdd.n740 iovdd.n738 0.818682
R762 iovdd.n930 iovdd.n929 0.818682
R763 iovdd.n928 iovdd.n927 0.818682
R764 iovdd.n746 iovdd.n745 0.818682
R765 iovdd.n920 iovdd.n919 0.818682
R766 iovdd.n918 iovdd.n917 0.818682
R767 iovdd.n810 iovdd.n809 0.818682
R768 iovdd.n818 iovdd.n816 0.818682
R769 iovdd.n909 iovdd.n908 0.818682
R770 iovdd.n907 iovdd.n906 0.818682
R771 iovdd.n824 iovdd.n823 0.818682
R772 iovdd.n831 iovdd.n829 0.818682
R773 iovdd.n898 iovdd.n897 0.818682
R774 iovdd.n896 iovdd.n895 0.818682
R775 iovdd.n837 iovdd.n836 0.818682
R776 iovdd.n843 iovdd.n841 0.818682
R777 iovdd.n887 iovdd.n886 0.818682
R778 iovdd.n885 iovdd.n884 0.818682
R779 iovdd.n849 iovdd.n848 0.818682
R780 iovdd.n857 iovdd.n855 0.818682
R781 iovdd.n876 iovdd.n875 0.818682
R782 iovdd.n874 iovdd.n873 0.818682
R783 iovdd.n863 iovdd.n862 0.818682
R784 iovdd.n1107 iovdd.n1106 0.818682
R785 iovdd.n5 iovdd.n4 0.818682
R786 iovdd.n1095 iovdd.n1094 0.818682
R787 iovdd.n1093 iovdd.n12 0.818682
R788 iovdd.n1092 iovdd.n1091 0.818682
R789 iovdd.n14 iovdd.n13 0.818682
R790 iovdd.n1079 iovdd.n1078 0.818682
R791 iovdd.n1077 iovdd.n23 0.818682
R792 iovdd.n1076 iovdd.n1075 0.818682
R793 iovdd.n25 iovdd.n24 0.818682
R794 iovdd.n1064 iovdd.n1063 0.818682
R795 iovdd.n1062 iovdd.n32 0.818682
R796 iovdd.n1061 iovdd.n1060 0.818682
R797 iovdd.n34 iovdd.n33 0.818682
R798 iovdd.n1049 iovdd.n1048 0.818682
R799 iovdd.n1047 iovdd.n41 0.818682
R800 iovdd.n1046 iovdd.n1045 0.818682
R801 iovdd.n43 iovdd.n42 0.818682
R802 iovdd.n1033 iovdd.n1032 0.818682
R803 iovdd.n1031 iovdd.n52 0.818682
R804 iovdd.n1030 iovdd.n1029 0.818682
R805 iovdd.n54 iovdd.n53 0.818682
R806 iovdd.n1018 iovdd.n1017 0.818682
R807 iovdd.n1016 iovdd.n61 0.818682
R808 iovdd.n1015 iovdd.n1014 0.818682
R809 iovdd.n63 iovdd.n62 0.818682
R810 iovdd.n1003 iovdd.n1002 0.818682
R811 iovdd.n1001 iovdd.n70 0.818682
R812 iovdd.n1000 iovdd.n999 0.818682
R813 iovdd.n72 iovdd.n71 0.818682
R814 iovdd.n987 iovdd.n986 0.818682
R815 iovdd.n985 iovdd.n961 0.818682
R816 iovdd.n984 iovdd.n983 0.818682
R817 iovdd.n963 iovdd.n962 0.818682
R818 iovdd.n972 iovdd.n971 0.818682
R819 iovdd.n969 iovdd.n967 0.818682
R820 iovdd.n973 iovdd.n972 0.818682
R821 iovdd.n964 iovdd.n963 0.818682
R822 iovdd.n983 iovdd.n982 0.818682
R823 iovdd.n961 iovdd.n959 0.818682
R824 iovdd.n988 iovdd.n987 0.818682
R825 iovdd.n73 iovdd.n72 0.818682
R826 iovdd.n999 iovdd.n998 0.818682
R827 iovdd.n70 iovdd.n68 0.818682
R828 iovdd.n1004 iovdd.n1003 0.818682
R829 iovdd.n64 iovdd.n63 0.818682
R830 iovdd.n1014 iovdd.n1013 0.818682
R831 iovdd.n61 iovdd.n59 0.818682
R832 iovdd.n1019 iovdd.n1018 0.818682
R833 iovdd.n55 iovdd.n54 0.818682
R834 iovdd.n1029 iovdd.n1028 0.818682
R835 iovdd.n52 iovdd.n50 0.818682
R836 iovdd.n1034 iovdd.n1033 0.818682
R837 iovdd.n44 iovdd.n43 0.818682
R838 iovdd.n1045 iovdd.n1044 0.818682
R839 iovdd.n41 iovdd.n39 0.818682
R840 iovdd.n1050 iovdd.n1049 0.818682
R841 iovdd.n35 iovdd.n34 0.818682
R842 iovdd.n1060 iovdd.n1059 0.818682
R843 iovdd.n32 iovdd.n30 0.818682
R844 iovdd.n1065 iovdd.n1064 0.818682
R845 iovdd.n26 iovdd.n25 0.818682
R846 iovdd.n1075 iovdd.n1074 0.818682
R847 iovdd.n23 iovdd.n21 0.818682
R848 iovdd.n1080 iovdd.n1079 0.818682
R849 iovdd.n15 iovdd.n14 0.818682
R850 iovdd.n1091 iovdd.n1090 0.818682
R851 iovdd.n12 iovdd.n10 0.818682
R852 iovdd.n1096 iovdd.n1095 0.818682
R853 iovdd.n6 iovdd.n5 0.818682
R854 iovdd.n1106 iovdd.n1105 0.818682
R855 iovdd.n3 iovdd.n2 0.818682
R856 iovdd.n626 iovdd.n625 0.762052
R857 iovdd.n603 iovdd.n602 0.698729
R858 iovdd.n602 iovdd.n601 0.698729
R859 iovdd.n601 iovdd.n600 0.698729
R860 iovdd.n401 iovdd.n400 0.698729
R861 iovdd.n402 iovdd.n401 0.698729
R862 iovdd.n403 iovdd.n402 0.698729
R863 iovdd.n392 iovdd.n391 0.698729
R864 iovdd.n393 iovdd.n392 0.698729
R865 iovdd.n394 iovdd.n393 0.698729
R866 iovdd.n378 iovdd.n377 0.698729
R867 iovdd.n379 iovdd.n378 0.698729
R868 iovdd.n380 iovdd.n379 0.698729
R869 iovdd.n368 iovdd.n367 0.698729
R870 iovdd.n369 iovdd.n368 0.698729
R871 iovdd.n370 iovdd.n369 0.698729
R872 iovdd.n354 iovdd.n353 0.698729
R873 iovdd.n355 iovdd.n354 0.698729
R874 iovdd.n356 iovdd.n355 0.698729
R875 iovdd.n344 iovdd.n343 0.698729
R876 iovdd.n345 iovdd.n344 0.698729
R877 iovdd.n346 iovdd.n345 0.698729
R878 iovdd.n331 iovdd.n330 0.698729
R879 iovdd.n332 iovdd.n331 0.698729
R880 iovdd.n333 iovdd.n332 0.698729
R881 iovdd.n314 iovdd.n313 0.698729
R882 iovdd.n315 iovdd.n314 0.698729
R883 iovdd.n316 iovdd.n315 0.698729
R884 iovdd.n306 iovdd.n305 0.698729
R885 iovdd.n307 iovdd.n306 0.698729
R886 iovdd.n308 iovdd.n307 0.698729
R887 iovdd.n297 iovdd.n296 0.698729
R888 iovdd.n298 iovdd.n297 0.698729
R889 iovdd.n299 iovdd.n298 0.698729
R890 iovdd.n283 iovdd.n282 0.698729
R891 iovdd.n284 iovdd.n283 0.698729
R892 iovdd.n285 iovdd.n284 0.698729
R893 iovdd.n273 iovdd.n272 0.698729
R894 iovdd.n274 iovdd.n273 0.698729
R895 iovdd.n275 iovdd.n274 0.698729
R896 iovdd.n259 iovdd.n258 0.698729
R897 iovdd.n260 iovdd.n259 0.698729
R898 iovdd.n261 iovdd.n260 0.698729
R899 iovdd.n249 iovdd.n248 0.698729
R900 iovdd.n250 iovdd.n249 0.698729
R901 iovdd.n251 iovdd.n250 0.698729
R902 iovdd.n236 iovdd.n235 0.698729
R903 iovdd.n237 iovdd.n236 0.698729
R904 iovdd.n238 iovdd.n237 0.698729
R905 iovdd.n221 iovdd.n220 0.698729
R906 iovdd.n222 iovdd.n221 0.698729
R907 iovdd.n223 iovdd.n222 0.698729
R908 iovdd.n212 iovdd.n211 0.698729
R909 iovdd.n213 iovdd.n212 0.698729
R910 iovdd.n214 iovdd.n213 0.698729
R911 iovdd.n205 iovdd.n204 0.698729
R912 iovdd.n206 iovdd.n205 0.698729
R913 iovdd.n207 iovdd.n206 0.698729
R914 iovdd.n160 iovdd.n159 0.698729
R915 iovdd.n161 iovdd.n160 0.698729
R916 iovdd.n162 iovdd.n161 0.698729
R917 iovdd.n169 iovdd.n168 0.698729
R918 iovdd.n170 iovdd.n169 0.698729
R919 iovdd.n171 iovdd.n170 0.698729
R920 iovdd.n610 iovdd.n609 0.698729
R921 iovdd.n611 iovdd.n610 0.698729
R922 iovdd.n612 iovdd.n611 0.698729
R923 iovdd.n608 iovdd.n607 0.564577
R924 iovdd.n659 iovdd.n46 0.548016
R925 iovdd.n656 iovdd.n46 0.548016
R926 iovdd.n653 iovdd.n46 0.548016
R927 iovdd.n650 iovdd.n46 0.548016
R928 iovdd.n642 iovdd.n18 0.548016
R929 iovdd.n639 iovdd.n18 0.548016
R930 iovdd.n636 iovdd.n18 0.548016
R931 iovdd.n633 iovdd.n18 0.548016
R932 iovdd.n607 iovdd.n116 0.526877
R933 iovdd.n605 iovdd.n604 0.496411
R934 iovdd.n605 iovdd.n139 0.471452
R935 iovdd.n700 iovdd.n690 0.416993
R936 iovdd.n971 iovdd.n970 0.416993
R937 iovdd.n1108 iovdd.n1107 0.416993
R938 iovdd.n761 iovdd.n760 0.328961
R939 iovdd.n795 iovdd.n794 0.328961
R940 iovdd.n599 iovdd.n140 0.323766
R941 iovdd.n774 iovdd.n773 0.322808
R942 iovdd.n783 iovdd.n782 0.322188
R943 iovdd.n600 iovdd 0.317156
R944 iovdd iovdd.n403 0.317156
R945 iovdd iovdd.n394 0.317156
R946 iovdd iovdd.n380 0.317156
R947 iovdd iovdd.n370 0.317156
R948 iovdd iovdd.n356 0.317156
R949 iovdd iovdd.n346 0.317156
R950 iovdd iovdd.n333 0.317156
R951 iovdd iovdd.n316 0.317156
R952 iovdd iovdd.n308 0.317156
R953 iovdd iovdd.n299 0.317156
R954 iovdd iovdd.n285 0.317156
R955 iovdd iovdd.n275 0.317156
R956 iovdd iovdd.n261 0.317156
R957 iovdd iovdd.n251 0.317156
R958 iovdd iovdd.n238 0.317156
R959 iovdd iovdd.n223 0.317156
R960 iovdd iovdd.n214 0.317156
R961 iovdd iovdd.n207 0.317156
R962 iovdd iovdd.n162 0.317156
R963 iovdd iovdd.n171 0.317156
R964 iovdd iovdd.n612 0.317156
R965 iovdd.n786 iovdd.n785 0.316029
R966 iovdd.n771 iovdd.n770 0.31602
R967 iovdd.n798 iovdd.n797 0.309867
R968 iovdd.n764 iovdd.n763 0.309867
R969 iovdd.n793 iovdd.n792 0.309247
R970 iovdd.n759 iovdd.n758 0.309247
R971 iovdd.n776 iovdd.n775 0.303088
R972 iovdd.n781 iovdd.n780 0.303079
R973 iovdd.n788 iovdd.n787 0.296926
R974 iovdd.n754 iovdd.n753 0.296926
R975 iovdd.n803 iovdd.n801 0.296305
R976 iovdd.n769 iovdd.n768 0.296305
R977 iovdd.n763 iovdd.n762 0.291089
R978 iovdd.n797 iovdd.n796 0.291089
R979 iovdd.n800 iovdd.n799 0.290146
R980 iovdd.n766 iovdd.n765 0.290146
R981 iovdd.n757 iovdd.n756 0.290137
R982 iovdd.n791 iovdd.n790 0.290137
R983 iovdd.n772 iovdd.n771 0.284975
R984 iovdd.n785 iovdd.n784 0.284443
R985 iovdd.n778 iovdd.n777 0.283985
R986 iovdd.n779 iovdd.n778 0.283364
R987 iovdd.n784 iovdd.n783 0.278673
R988 iovdd.n773 iovdd.n772 0.278148
R989 iovdd.n790 iovdd.n789 0.277205
R990 iovdd.n756 iovdd.n755 0.277205
R991 iovdd.n767 iovdd.n766 0.277196
R992 iovdd.n802 iovdd.n800 0.277196
R993 iovdd.n762 iovdd.n761 0.272034
R994 iovdd.n796 iovdd.n795 0.272034
R995 iovdd.n803 iovdd.n802 0.271044
R996 iovdd.n768 iovdd.n767 0.271044
R997 iovdd.n789 iovdd.n788 0.270423
R998 iovdd.n755 iovdd.n754 0.270423
R999 iovdd.n780 iovdd.n779 0.264264
R1000 iovdd.n777 iovdd.n776 0.264255
R1001 iovdd.n329 iovdd.n130 0.262329
R1002 iovdd.n399 iovdd.n115 0.259848
R1003 iovdd.n203 iovdd.n120 0.259729
R1004 iovdd.n234 iovdd.n122 0.258965
R1005 iovdd.n792 iovdd.n791 0.258102
R1006 iovdd.n758 iovdd.n757 0.258102
R1007 iovdd.n799 iovdd.n798 0.257482
R1008 iovdd.n765 iovdd.n764 0.257482
R1009 iovdd.n295 iovdd.n128 0.256612
R1010 iovdd.n342 iovdd.n131 0.255729
R1011 iovdd.n158 iovdd.n119 0.253377
R1012 iovdd.n390 iovdd.n136 0.253259
R1013 iovdd.n247 iovdd.n123 0.252623
R1014 iovdd.n770 iovdd.n769 0.251323
R1015 iovdd.n787 iovdd.n786 0.251314
R1016 iovdd.n281 iovdd.n127 0.250024
R1017 iovdd.n352 iovdd.n132 0.249388
R1018 iovdd.n149 iovdd 0.248
R1019 iovdd.n376 iovdd.n135 0.246906
R1020 iovdd.n167 iovdd.n118 0.246788
R1021 iovdd.n257 iovdd.n124 0.246024
R1022 iovdd.n782 iovdd.n781 0.245161
R1023 iovdd.n775 iovdd.n774 0.244541
R1024 iovdd.n312 iovdd.n129 0.243764
R1025 iovdd.n271 iovdd.n126 0.243671
R1026 iovdd.n366 iovdd.n133 0.242788
R1027 iovdd.n210 iovdd.n121 0.241516
R1028 iovdd.n606 iovdd.n605 0.241185
R1029 iovdd.n604 iovdd.n117 0.240436
R1030 iovdd.n366 iovdd.n134 0.240318
R1031 iovdd.n219 iovdd.n121 0.24031
R1032 iovdd.n271 iovdd.n125 0.239682
R1033 iovdd.n794 iovdd.n793 0.238382
R1034 iovdd.n760 iovdd.n759 0.238382
R1035 iovdd.n304 iovdd.n129 0.238095
R1036 iovdd.n257 iovdd.n125 0.237082
R1037 iovdd.n376 iovdd.n134 0.236447
R1038 iovdd.n167 iovdd.n117 0.236318
R1039 iovdd.n352 iovdd.n133 0.233965
R1040 iovdd.n281 iovdd.n126 0.233082
R1041 iovdd.n247 iovdd.n124 0.23073
R1042 iovdd.n158 iovdd.n118 0.229976
R1043 iovdd.n390 iovdd.n135 0.229847
R1044 iovdd.n342 iovdd.n132 0.227377
R1045 iovdd.n295 iovdd.n127 0.226741
R1046 iovdd.n234 iovdd.n123 0.224141
R1047 iovdd.n399 iovdd.n136 0.223506
R1048 iovdd.n203 iovdd.n119 0.223377
R1049 iovdd.n329 iovdd.n131 0.221024
R1050 iovdd.n304 iovdd.n128 0.220141
R1051 iovdd.n219 iovdd.n122 0.217789
R1052 iovdd.n210 iovdd.n120 0.217035
R1053 iovdd.n608 iovdd.n115 0.216906
R1054 iovdd.n312 iovdd.n130 0.214435
R1055 iovdd.n694 iovdd.n693 0.201704
R1056 iovdd.n976 iovdd.n966 0.201704
R1057 iovdd.n868 iovdd.n867 0.2005
R1058 iovdd.n872 iovdd.n871 0.2005
R1059 iovdd.n856 iovdd.n853 0.2005
R1060 iovdd.n878 iovdd.n877 0.2005
R1061 iovdd.n854 iovdd.n850 0.2005
R1062 iovdd.n883 iovdd.n882 0.2005
R1063 iovdd.n842 iovdd.n839 0.2005
R1064 iovdd.n889 iovdd.n888 0.2005
R1065 iovdd.n840 iovdd.n838 0.2005
R1066 iovdd.n894 iovdd.n893 0.2005
R1067 iovdd.n830 iovdd.n827 0.2005
R1068 iovdd.n900 iovdd.n899 0.2005
R1069 iovdd.n828 iovdd.n825 0.2005
R1070 iovdd.n905 iovdd.n904 0.2005
R1071 iovdd.n817 iovdd.n814 0.2005
R1072 iovdd.n911 iovdd.n910 0.2005
R1073 iovdd.n815 iovdd.n811 0.2005
R1074 iovdd.n916 iovdd.n915 0.2005
R1075 iovdd.n748 iovdd.n747 0.2005
R1076 iovdd.n922 iovdd.n921 0.2005
R1077 iovdd.n926 iovdd.n925 0.2005
R1078 iovdd.n739 iovdd.n736 0.2005
R1079 iovdd.n932 iovdd.n931 0.2005
R1080 iovdd.n737 iovdd.n734 0.2005
R1081 iovdd.n937 iovdd.n936 0.2005
R1082 iovdd.n726 iovdd.n723 0.2005
R1083 iovdd.n943 iovdd.n942 0.2005
R1084 iovdd.n724 iovdd.n721 0.2005
R1085 iovdd.n948 iovdd.n947 0.2005
R1086 iovdd.n679 iovdd.n677 0.2005
R1087 iovdd.n954 iovdd.n953 0.2005
R1088 iovdd.n712 iovdd.n676 0.2005
R1089 iovdd.n711 iovdd.n710 0.2005
R1090 iovdd.n688 iovdd.n684 0.2005
R1091 iovdd.n706 iovdd.n705 0.2005
R1092 iovdd.n697 iovdd.n686 0.2005
R1093 iovdd.n696 iovdd.n695 0.2005
R1094 iovdd.n1110 iovdd.n1109 0.2005
R1095 iovdd.n1104 iovdd.n1 0.2005
R1096 iovdd.n1103 iovdd.n1102 0.2005
R1097 iovdd.n11 iovdd.n7 0.2005
R1098 iovdd.n1098 iovdd.n1097 0.2005
R1099 iovdd.n1089 iovdd.n9 0.2005
R1100 iovdd.n1088 iovdd.n1087 0.2005
R1101 iovdd.n22 iovdd.n16 0.2005
R1102 iovdd.n1082 iovdd.n1081 0.2005
R1103 iovdd.n1073 iovdd.n20 0.2005
R1104 iovdd.n1072 iovdd.n1071 0.2005
R1105 iovdd.n31 iovdd.n27 0.2005
R1106 iovdd.n1067 iovdd.n1066 0.2005
R1107 iovdd.n1058 iovdd.n29 0.2005
R1108 iovdd.n1057 iovdd.n1056 0.2005
R1109 iovdd.n40 iovdd.n36 0.2005
R1110 iovdd.n1052 iovdd.n1051 0.2005
R1111 iovdd.n1043 iovdd.n38 0.2005
R1112 iovdd.n1042 iovdd.n1041 0.2005
R1113 iovdd.n51 iovdd.n45 0.2005
R1114 iovdd.n1036 iovdd.n1035 0.2005
R1115 iovdd.n1027 iovdd.n49 0.2005
R1116 iovdd.n1026 iovdd.n1025 0.2005
R1117 iovdd.n60 iovdd.n56 0.2005
R1118 iovdd.n1021 iovdd.n1020 0.2005
R1119 iovdd.n1012 iovdd.n58 0.2005
R1120 iovdd.n1011 iovdd.n1010 0.2005
R1121 iovdd.n69 iovdd.n65 0.2005
R1122 iovdd.n1006 iovdd.n1005 0.2005
R1123 iovdd.n997 iovdd.n67 0.2005
R1124 iovdd.n996 iovdd.n995 0.2005
R1125 iovdd.n960 iovdd.n74 0.2005
R1126 iovdd.n990 iovdd.n989 0.2005
R1127 iovdd.n981 iovdd.n958 0.2005
R1128 iovdd.n980 iovdd.n979 0.2005
R1129 iovdd.n968 iovdd.n965 0.2005
R1130 iovdd.n975 iovdd.n974 0.2005
R1131 iovdd.n607 iovdd.n606 0.173189
R1132 iovdd.n804 iovdd.n752 0.166751
R1133 iovdd.n46 iovdd 0.16242
R1134 iovdd.n807 iovdd.n806 0.156347
R1135 iovdd.n109 iovdd 0.119054
R1136 iovdd.n869 iovdd.n868 0.1105
R1137 iovdd.n871 iovdd.n870 0.1105
R1138 iovdd.n853 iovdd.n852 0.1105
R1139 iovdd.n879 iovdd.n878 0.1105
R1140 iovdd.n880 iovdd.n850 0.1105
R1141 iovdd.n882 iovdd.n881 0.1105
R1142 iovdd.n851 iovdd.n839 0.1105
R1143 iovdd.n890 iovdd.n889 0.1105
R1144 iovdd.n891 iovdd.n838 0.1105
R1145 iovdd.n893 iovdd.n892 0.1105
R1146 iovdd.n827 iovdd.n826 0.1105
R1147 iovdd.n901 iovdd.n900 0.1105
R1148 iovdd.n902 iovdd.n825 0.1105
R1149 iovdd.n904 iovdd.n903 0.1105
R1150 iovdd.n814 iovdd.n813 0.1105
R1151 iovdd.n912 iovdd.n911 0.1105
R1152 iovdd.n913 iovdd.n811 0.1105
R1153 iovdd.n915 iovdd.n914 0.1105
R1154 iovdd.n812 iovdd.n747 0.1105
R1155 iovdd.n923 iovdd.n922 0.1105
R1156 iovdd.n925 iovdd.n924 0.1105
R1157 iovdd.n736 iovdd.n735 0.1105
R1158 iovdd.n933 iovdd.n932 0.1105
R1159 iovdd.n934 iovdd.n734 0.1105
R1160 iovdd.n936 iovdd.n935 0.1105
R1161 iovdd.n723 iovdd.n722 0.1105
R1162 iovdd.n944 iovdd.n943 0.1105
R1163 iovdd.n945 iovdd.n721 0.1105
R1164 iovdd.n947 iovdd.n946 0.1105
R1165 iovdd.n677 iovdd.n675 0.1105
R1166 iovdd.n955 iovdd.n954 0.1105
R1167 iovdd.n676 iovdd.n674 0.1105
R1168 iovdd.n710 iovdd.n709 0.1105
R1169 iovdd.n708 iovdd.n684 0.1105
R1170 iovdd.n707 iovdd.n706 0.1105
R1171 iovdd.n686 iovdd.n685 0.1105
R1172 iovdd.n1111 iovdd.n1110 0.1105
R1173 iovdd.n1 iovdd.n0 0.1105
R1174 iovdd.n1102 iovdd.n1101 0.1105
R1175 iovdd.n1100 iovdd.n7 0.1105
R1176 iovdd.n1099 iovdd.n1098 0.1105
R1177 iovdd.n9 iovdd.n8 0.1105
R1178 iovdd.n1087 iovdd.n1086 0.1105
R1179 iovdd.n1084 iovdd.n16 0.1105
R1180 iovdd.n1083 iovdd.n1082 0.1105
R1181 iovdd.n20 iovdd.n19 0.1105
R1182 iovdd.n1071 iovdd.n1070 0.1105
R1183 iovdd.n1069 iovdd.n27 0.1105
R1184 iovdd.n1068 iovdd.n1067 0.1105
R1185 iovdd.n29 iovdd.n28 0.1105
R1186 iovdd.n1056 iovdd.n1055 0.1105
R1187 iovdd.n1054 iovdd.n36 0.1105
R1188 iovdd.n1053 iovdd.n1052 0.1105
R1189 iovdd.n38 iovdd.n37 0.1105
R1190 iovdd.n1041 iovdd.n1040 0.1105
R1191 iovdd.n1038 iovdd.n45 0.1105
R1192 iovdd.n1037 iovdd.n1036 0.1105
R1193 iovdd.n49 iovdd.n48 0.1105
R1194 iovdd.n1025 iovdd.n1024 0.1105
R1195 iovdd.n1023 iovdd.n56 0.1105
R1196 iovdd.n1022 iovdd.n1021 0.1105
R1197 iovdd.n58 iovdd.n57 0.1105
R1198 iovdd.n1010 iovdd.n1009 0.1105
R1199 iovdd.n1008 iovdd.n65 0.1105
R1200 iovdd.n1007 iovdd.n1006 0.1105
R1201 iovdd.n67 iovdd.n66 0.1105
R1202 iovdd.n995 iovdd.n994 0.1105
R1203 iovdd.n992 iovdd.n74 0.1105
R1204 iovdd.n991 iovdd.n990 0.1105
R1205 iovdd.n958 iovdd.n957 0.1105
R1206 iovdd.n979 iovdd.n978 0.1105
R1207 iovdd.n977 iovdd.n965 0.1105
R1208 iovdd.n18 iovdd 0.0768767
R1209 iovdd.n595 iovdd.n143 0.0591667
R1210 iovdd.n595 iovdd.n144 0.0591667
R1211 iovdd.n184 iovdd.n144 0.0591667
R1212 iovdd.n184 iovdd.n152 0.0591667
R1213 iovdd.n585 iovdd.n152 0.0591667
R1214 iovdd.n585 iovdd.n153 0.0591667
R1215 iovdd.n229 iovdd.n153 0.0591667
R1216 iovdd.n230 iovdd.n229 0.0591667
R1217 iovdd.n554 iovdd.n230 0.0591667
R1218 iovdd.n554 iovdd.n552 0.0591667
R1219 iovdd.n552 iovdd.n231 0.0591667
R1220 iovdd.n535 iovdd.n231 0.0591667
R1221 iovdd.n535 iovdd.n534 0.0591667
R1222 iovdd.n534 iovdd.n254 0.0591667
R1223 iovdd.n517 iovdd.n254 0.0591667
R1224 iovdd.n517 iovdd.n516 0.0591667
R1225 iovdd.n516 iovdd.n278 0.0591667
R1226 iovdd.n322 iovdd.n278 0.0591667
R1227 iovdd.n323 iovdd.n322 0.0591667
R1228 iovdd.n324 iovdd.n323 0.0591667
R1229 iovdd.n478 iovdd.n324 0.0591667
R1230 iovdd.n478 iovdd.n477 0.0591667
R1231 iovdd.n477 iovdd.n326 0.0591667
R1232 iovdd.n460 iovdd.n326 0.0591667
R1233 iovdd.n460 iovdd.n459 0.0591667
R1234 iovdd.n459 iovdd.n349 0.0591667
R1235 iovdd.n442 iovdd.n349 0.0591667
R1236 iovdd.n442 iovdd.n441 0.0591667
R1237 iovdd.n441 iovdd.n373 0.0591667
R1238 iovdd.n406 iovdd.n373 0.0591667
R1239 iovdd.n407 iovdd.n406 0.0591667
R1240 iovdd.n408 iovdd.n407 0.0591667
R1241 iovdd.n408 iovdd.n107 0.0591667
R1242 iovdd.n627 iovdd.n107 0.0591667
R1243 iovdd.n594 iovdd.n145 0.0591667
R1244 iovdd.n594 iovdd.n146 0.0591667
R1245 iovdd.n151 iovdd.n146 0.0591667
R1246 iovdd.n587 iovdd.n151 0.0591667
R1247 iovdd.n587 iovdd.n586 0.0591667
R1248 iovdd.n586 iovdd.n78 0.0591667
R1249 iovdd.n79 iovdd.n78 0.0591667
R1250 iovdd.n80 iovdd.n79 0.0591667
R1251 iovdd.n553 iovdd.n80 0.0591667
R1252 iovdd.n553 iovdd.n83 0.0591667
R1253 iovdd.n84 iovdd.n83 0.0591667
R1254 iovdd.n85 iovdd.n84 0.0591667
R1255 iovdd.n86 iovdd.n85 0.0591667
R1256 iovdd.n87 iovdd.n86 0.0591667
R1257 iovdd.n88 iovdd.n87 0.0591667
R1258 iovdd.n89 iovdd.n88 0.0591667
R1259 iovdd.n90 iovdd.n89 0.0591667
R1260 iovdd.n91 iovdd.n90 0.0591667
R1261 iovdd.n92 iovdd.n91 0.0591667
R1262 iovdd.n93 iovdd.n92 0.0591667
R1263 iovdd.n94 iovdd.n93 0.0591667
R1264 iovdd.n95 iovdd.n94 0.0591667
R1265 iovdd.n325 iovdd.n95 0.0591667
R1266 iovdd.n325 iovdd.n97 0.0591667
R1267 iovdd.n98 iovdd.n97 0.0591667
R1268 iovdd.n99 iovdd.n98 0.0591667
R1269 iovdd.n100 iovdd.n99 0.0591667
R1270 iovdd.n101 iovdd.n100 0.0591667
R1271 iovdd.n102 iovdd.n101 0.0591667
R1272 iovdd.n103 iovdd.n102 0.0591667
R1273 iovdd.n104 iovdd.n103 0.0591667
R1274 iovdd.n105 iovdd.n104 0.0591667
R1275 iovdd.n106 iovdd.n105 0.0591667
R1276 iovdd.n628 iovdd.n106 0.0591667
R1277 iovdd.n694 iovdd.n685 0.0568704
R1278 iovdd.n977 iovdd.n976 0.0568704
R1279 iovdd.n751 iovdd 0.0555
R1280 iovdd.n804 iovdd.t89 0.0507959
R1281 iovdd.n1039 iovdd.n46 0.0401072
R1282 iovdd.n1085 iovdd.n18 0.0401072
R1283 iovdd.n597 iovdd.n140 0.0374917
R1284 iovdd.n625 iovdd.n624 0.02024
R1285 iovdd.n598 iovdd.n141 0.0148733
R1286 iovdd.n173 iovdd.n141 0.0148733
R1287 iovdd.n173 iovdd.n172 0.0148733
R1288 iovdd.n178 iovdd.n172 0.0148733
R1289 iovdd.n179 iovdd.n178 0.0148733
R1290 iovdd.n181 iovdd.n165 0.0148733
R1291 iovdd.n187 iovdd.n165 0.0148733
R1292 iovdd.n188 iovdd.n187 0.0148733
R1293 iovdd.n189 iovdd.n188 0.0148733
R1294 iovdd.n189 iovdd.n163 0.0148733
R1295 iovdd.n194 iovdd.n163 0.0148733
R1296 iovdd.n197 iovdd.n196 0.0148733
R1297 iovdd.n197 iovdd.n156 0.0148733
R1298 iovdd.n201 iovdd.n156 0.0148733
R1299 iovdd.n202 iovdd.n201 0.0148733
R1300 iovdd.n582 iovdd.n202 0.0148733
R1301 iovdd.n580 iovdd.n579 0.0148733
R1302 iovdd.n579 iovdd.n208 0.0148733
R1303 iovdd.n574 iovdd.n208 0.0148733
R1304 iovdd.n574 iovdd.n573 0.0148733
R1305 iovdd.n573 iovdd.n572 0.0148733
R1306 iovdd.n569 iovdd.n568 0.0148733
R1307 iovdd.n568 iovdd.n217 0.0148733
R1308 iovdd.n564 iovdd.n217 0.0148733
R1309 iovdd.n564 iovdd.n563 0.0148733
R1310 iovdd.n563 iovdd.n562 0.0148733
R1311 iovdd.n559 iovdd.n558 0.0148733
R1312 iovdd.n558 iovdd.n557 0.0148733
R1313 iovdd.n557 iovdd.n227 0.0148733
R1314 iovdd.n239 iovdd.n227 0.0148733
R1315 iovdd.n242 iovdd.n239 0.0148733
R1316 iovdd.n549 iovdd.n244 0.0148733
R1317 iovdd.n549 iovdd.n548 0.0148733
R1318 iovdd.n548 iovdd.n547 0.0148733
R1319 iovdd.n547 iovdd.n245 0.0148733
R1320 iovdd.n542 iovdd.n245 0.0148733
R1321 iovdd.n540 iovdd.n539 0.0148733
R1322 iovdd.n539 iovdd.n252 0.0148733
R1323 iovdd.n262 iovdd.n252 0.0148733
R1324 iovdd.n263 iovdd.n262 0.0148733
R1325 iovdd.n266 iovdd.n263 0.0148733
R1326 iovdd.n267 iovdd.n266 0.0148733
R1327 iovdd.n531 iovdd.n530 0.0148733
R1328 iovdd.n530 iovdd.n529 0.0148733
R1329 iovdd.n529 iovdd.n269 0.0148733
R1330 iovdd.n524 iovdd.n269 0.0148733
R1331 iovdd.n524 iovdd.n523 0.0148733
R1332 iovdd.n521 iovdd.n276 0.0148733
R1333 iovdd.n286 iovdd.n276 0.0148733
R1334 iovdd.n287 iovdd.n286 0.0148733
R1335 iovdd.n290 iovdd.n287 0.0148733
R1336 iovdd.n291 iovdd.n290 0.0148733
R1337 iovdd.n513 iovdd.n512 0.0148733
R1338 iovdd.n512 iovdd.n511 0.0148733
R1339 iovdd.n511 iovdd.n293 0.0148733
R1340 iovdd.n507 iovdd.n293 0.0148733
R1341 iovdd.n507 iovdd.n506 0.0148733
R1342 iovdd.n504 iovdd.n300 0.0148733
R1343 iovdd.n500 iovdd.n300 0.0148733
R1344 iovdd.n500 iovdd.n499 0.0148733
R1345 iovdd.n499 iovdd.n302 0.0148733
R1346 iovdd.n495 iovdd.n302 0.0148733
R1347 iovdd.n493 iovdd.n492 0.0148733
R1348 iovdd.n492 iovdd.n309 0.0148733
R1349 iovdd.n488 iovdd.n309 0.0148733
R1350 iovdd.n488 iovdd.n487 0.0148733
R1351 iovdd.n487 iovdd.n486 0.0148733
R1352 iovdd.n483 iovdd.n482 0.0148733
R1353 iovdd.n482 iovdd.n481 0.0148733
R1354 iovdd.n481 iovdd.n320 0.0148733
R1355 iovdd.n334 iovdd.n320 0.0148733
R1356 iovdd.n337 iovdd.n334 0.0148733
R1357 iovdd.n338 iovdd.n337 0.0148733
R1358 iovdd.n474 iovdd.n473 0.0148733
R1359 iovdd.n473 iovdd.n472 0.0148733
R1360 iovdd.n472 iovdd.n340 0.0148733
R1361 iovdd.n467 iovdd.n340 0.0148733
R1362 iovdd.n467 iovdd.n466 0.0148733
R1363 iovdd.n464 iovdd.n347 0.0148733
R1364 iovdd.n357 iovdd.n347 0.0148733
R1365 iovdd.n358 iovdd.n357 0.0148733
R1366 iovdd.n361 iovdd.n358 0.0148733
R1367 iovdd.n362 iovdd.n361 0.0148733
R1368 iovdd.n456 iovdd.n455 0.0148733
R1369 iovdd.n455 iovdd.n454 0.0148733
R1370 iovdd.n454 iovdd.n364 0.0148733
R1371 iovdd.n449 iovdd.n364 0.0148733
R1372 iovdd.n449 iovdd.n448 0.0148733
R1373 iovdd.n446 iovdd.n371 0.0148733
R1374 iovdd.n381 iovdd.n371 0.0148733
R1375 iovdd.n382 iovdd.n381 0.0148733
R1376 iovdd.n385 iovdd.n382 0.0148733
R1377 iovdd.n386 iovdd.n385 0.0148733
R1378 iovdd.n438 iovdd.n437 0.0148733
R1379 iovdd.n437 iovdd.n436 0.0148733
R1380 iovdd.n436 iovdd.n388 0.0148733
R1381 iovdd.n431 iovdd.n388 0.0148733
R1382 iovdd.n431 iovdd.n430 0.0148733
R1383 iovdd.n428 iovdd.n395 0.0148733
R1384 iovdd.n424 iovdd.n395 0.0148733
R1385 iovdd.n424 iovdd.n423 0.0148733
R1386 iovdd.n423 iovdd.n397 0.0148733
R1387 iovdd.n419 iovdd.n397 0.0148733
R1388 iovdd.n419 iovdd.n418 0.0148733
R1389 iovdd.n416 iovdd.n404 0.0148733
R1390 iovdd.n412 iovdd.n404 0.0148733
R1391 iovdd.n412 iovdd.n411 0.0148733
R1392 iovdd.n411 iovdd.n114 0.0148733
R1393 iovdd.n614 iovdd.n114 0.0148733
R1394 iovdd.n618 iovdd.n112 0.0148733
R1395 iovdd.n619 iovdd.n618 0.0148733
R1396 iovdd.n619 iovdd.n110 0.0148733
R1397 iovdd.n623 iovdd.n110 0.0148733
R1398 iovdd.n624 iovdd.n623 0.0148733
R1399 iovdd.n174 iovdd.n142 0.0148733
R1400 iovdd.n175 iovdd.n174 0.0148733
R1401 iovdd.n177 iovdd.n175 0.0148733
R1402 iovdd.n182 iovdd.n166 0.0148733
R1403 iovdd.n183 iovdd.n182 0.0148733
R1404 iovdd.n186 iovdd.n183 0.0148733
R1405 iovdd.n190 iovdd.n164 0.0148733
R1406 iovdd.n191 iovdd.n190 0.0148733
R1407 iovdd.n193 iovdd.n191 0.0148733
R1408 iovdd.n198 iovdd.n157 0.0148733
R1409 iovdd.n199 iovdd.n198 0.0148733
R1410 iovdd.n200 iovdd.n199 0.0148733
R1411 iovdd.n200 iovdd.n154 0.0148733
R1412 iovdd.n583 iovdd.n155 0.0148733
R1413 iovdd.n578 iovdd.n155 0.0148733
R1414 iovdd.n578 iovdd.n577 0.0148733
R1415 iovdd.n575 iovdd.n209 0.0148733
R1416 iovdd.n571 iovdd.n209 0.0148733
R1417 iovdd.n571 iovdd.n570 0.0148733
R1418 iovdd.n567 iovdd.n566 0.0148733
R1419 iovdd.n566 iovdd.n565 0.0148733
R1420 iovdd.n565 iovdd.n218 0.0148733
R1421 iovdd.n561 iovdd.n560 0.0148733
R1422 iovdd.n560 iovdd.n226 0.0148733
R1423 iovdd.n556 iovdd.n226 0.0148733
R1424 iovdd.n240 iovdd.n228 0.0148733
R1425 iovdd.n241 iovdd.n240 0.0148733
R1426 iovdd.n241 iovdd.n232 0.0148733
R1427 iovdd.n550 iovdd.n233 0.0148733
R1428 iovdd.n546 iovdd.n233 0.0148733
R1429 iovdd.n546 iovdd.n545 0.0148733
R1430 iovdd.n543 iovdd.n246 0.0148733
R1431 iovdd.n538 iovdd.n246 0.0148733
R1432 iovdd.n538 iovdd.n537 0.0148733
R1433 iovdd.n264 iovdd.n253 0.0148733
R1434 iovdd.n265 iovdd.n264 0.0148733
R1435 iovdd.n265 iovdd.n255 0.0148733
R1436 iovdd.n532 iovdd.n256 0.0148733
R1437 iovdd.n528 iovdd.n256 0.0148733
R1438 iovdd.n528 iovdd.n527 0.0148733
R1439 iovdd.n525 iovdd.n270 0.0148733
R1440 iovdd.n520 iovdd.n270 0.0148733
R1441 iovdd.n520 iovdd.n519 0.0148733
R1442 iovdd.n288 iovdd.n277 0.0148733
R1443 iovdd.n289 iovdd.n288 0.0148733
R1444 iovdd.n289 iovdd.n279 0.0148733
R1445 iovdd.n514 iovdd.n280 0.0148733
R1446 iovdd.n510 iovdd.n280 0.0148733
R1447 iovdd.n510 iovdd.n509 0.0148733
R1448 iovdd.n509 iovdd.n508 0.0148733
R1449 iovdd.n508 iovdd.n294 0.0148733
R1450 iovdd.n503 iovdd.n294 0.0148733
R1451 iovdd.n503 iovdd.n502 0.0148733
R1452 iovdd.n502 iovdd.n501 0.0148733
R1453 iovdd.n498 iovdd.n497 0.0148733
R1454 iovdd.n497 iovdd.n496 0.0148733
R1455 iovdd.n496 iovdd.n303 0.0148733
R1456 iovdd.n491 iovdd.n490 0.0148733
R1457 iovdd.n490 iovdd.n489 0.0148733
R1458 iovdd.n489 iovdd.n311 0.0148733
R1459 iovdd.n485 iovdd.n484 0.0148733
R1460 iovdd.n484 iovdd.n319 0.0148733
R1461 iovdd.n480 iovdd.n319 0.0148733
R1462 iovdd.n335 iovdd.n321 0.0148733
R1463 iovdd.n336 iovdd.n335 0.0148733
R1464 iovdd.n336 iovdd.n327 0.0148733
R1465 iovdd.n475 iovdd.n328 0.0148733
R1466 iovdd.n471 iovdd.n328 0.0148733
R1467 iovdd.n471 iovdd.n470 0.0148733
R1468 iovdd.n468 iovdd.n341 0.0148733
R1469 iovdd.n463 iovdd.n341 0.0148733
R1470 iovdd.n463 iovdd.n462 0.0148733
R1471 iovdd.n359 iovdd.n348 0.0148733
R1472 iovdd.n360 iovdd.n359 0.0148733
R1473 iovdd.n360 iovdd.n350 0.0148733
R1474 iovdd.n457 iovdd.n351 0.0148733
R1475 iovdd.n453 iovdd.n351 0.0148733
R1476 iovdd.n453 iovdd.n452 0.0148733
R1477 iovdd.n450 iovdd.n365 0.0148733
R1478 iovdd.n445 iovdd.n365 0.0148733
R1479 iovdd.n445 iovdd.n444 0.0148733
R1480 iovdd.n383 iovdd.n372 0.0148733
R1481 iovdd.n384 iovdd.n383 0.0148733
R1482 iovdd.n384 iovdd.n374 0.0148733
R1483 iovdd.n439 iovdd.n375 0.0148733
R1484 iovdd.n435 iovdd.n375 0.0148733
R1485 iovdd.n435 iovdd.n434 0.0148733
R1486 iovdd.n432 iovdd.n389 0.0148733
R1487 iovdd.n427 iovdd.n389 0.0148733
R1488 iovdd.n427 iovdd.n426 0.0148733
R1489 iovdd.n426 iovdd.n425 0.0148733
R1490 iovdd.n422 iovdd.n421 0.0148733
R1491 iovdd.n421 iovdd.n420 0.0148733
R1492 iovdd.n420 iovdd.n398 0.0148733
R1493 iovdd.n415 iovdd.n414 0.0148733
R1494 iovdd.n414 iovdd.n413 0.0148733
R1495 iovdd.n413 iovdd.n410 0.0148733
R1496 iovdd.n615 iovdd.n113 0.0148733
R1497 iovdd.n616 iovdd.n615 0.0148733
R1498 iovdd.n617 iovdd.n616 0.0148733
R1499 iovdd.n621 iovdd.n620 0.0148733
R1500 iovdd.n622 iovdd.n621 0.0148733
R1501 iovdd.n622 iovdd.n108 0.0148733
R1502 iovdd.n417 iovdd.n416 0.0147267
R1503 iovdd.n584 iovdd.n583 0.01458
R1504 iovdd.n434 iovdd.n433 0.01458
R1505 iovdd.n474 iovdd.n339 0.0144333
R1506 iovdd.n805 iovdd.n804 0.0142662
R1507 iovdd.n531 iovdd.n268 0.01414
R1508 iovdd.n193 iovdd.n192 0.0139933
R1509 iovdd.n422 iovdd.n396 0.0139933
R1510 iovdd.n196 iovdd.n195 0.0138467
R1511 iovdd.n515 iovdd.n279 0.0137
R1512 iovdd.n498 iovdd.n301 0.0137
R1513 iovdd.n180 iovdd.n179 0.0135533
R1514 iovdd.n576 iovdd.n575 0.0134067
R1515 iovdd.n440 iovdd.n374 0.0134067
R1516 iovdd.n542 iovdd.n541 0.01326
R1517 iovdd.n486 iovdd.n317 0.0129667
R1518 iovdd.n186 iovdd.n185 0.01282
R1519 iovdd.n415 iovdd.n405 0.01282
R1520 iovdd.n430 iovdd.n429 0.0126733
R1521 iovdd.n519 iovdd.n518 0.0125267
R1522 iovdd.n491 iovdd.n310 0.0125267
R1523 iovdd.n593 iovdd.n147 0.0125
R1524 iovdd.n593 iovdd.n148 0.0125
R1525 iovdd.n589 iovdd.n148 0.0125
R1526 iovdd.n589 iovdd.n588 0.0125
R1527 iovdd.n588 iovdd.n77 0.0125
R1528 iovdd.n672 iovdd.n77 0.0125
R1529 iovdd.n672 iovdd.n671 0.0125
R1530 iovdd.n671 iovdd.n670 0.0125
R1531 iovdd.n670 iovdd.n81 0.0125
R1532 iovdd.n665 iovdd.n81 0.0125
R1533 iovdd.n665 iovdd.n664 0.0125
R1534 iovdd.n664 iovdd.n663 0.0125
R1535 iovdd.n663 iovdd.n661 0.0125
R1536 iovdd.n661 iovdd.n660 0.0125
R1537 iovdd.n658 iovdd.n657 0.0125
R1538 iovdd.n655 iovdd.n654 0.0125
R1539 iovdd.n652 iovdd.n651 0.0125
R1540 iovdd.n649 iovdd.n648 0.0125
R1541 iovdd.n648 iovdd.n96 0.0125
R1542 iovdd.n644 iovdd.n96 0.0125
R1543 iovdd.n644 iovdd.n643 0.0125
R1544 iovdd.n641 iovdd.n640 0.0125
R1545 iovdd.n638 iovdd.n637 0.0125
R1546 iovdd.n635 iovdd.n634 0.0125
R1547 iovdd.n632 iovdd.n631 0.0125
R1548 iovdd.n631 iovdd.n630 0.0125
R1549 iovdd.n613 iovdd.n112 0.01238
R1550 iovdd.n567 iovdd.n216 0.0122333
R1551 iovdd.n444 iovdd.n443 0.0122333
R1552 iovdd.n465 iovdd.n464 0.0120867
R1553 iovdd.n522 iovdd.n521 0.0117933
R1554 iovdd.n177 iovdd.n176 0.0116467
R1555 iovdd.n409 iovdd.n113 0.0116467
R1556 iovdd.n581 iovdd.n580 0.0115
R1557 iovdd.n527 iovdd.n526 0.0113533
R1558 iovdd.n485 iovdd.n318 0.0113533
R1559 iovdd.n561 iovdd.n225 0.01106
R1560 iovdd.n452 iovdd.n451 0.01106
R1561 iovdd.n243 iovdd.n242 0.0109133
R1562 iovdd.n495 iovdd.n494 0.01062
R1563 iovdd.n597 iovdd.n596 0.0104733
R1564 iovdd.n620 iovdd.n111 0.0104733
R1565 iovdd.n387 iovdd.n386 0.0103267
R1566 iovdd.n533 iovdd.n255 0.01018
R1567 iovdd.n479 iovdd.n321 0.01018
R1568 iovdd.n555 iovdd.n228 0.00988667
R1569 iovdd.n458 iovdd.n350 0.00988667
R1570 iovdd.n456 iovdd.n363 0.00974
R1571 iovdd.n513 iovdd.n292 0.00944667
R1572 iovdd.n569 iovdd.n215 0.00915333
R1573 iovdd.n537 iovdd.n536 0.00900667
R1574 iovdd.n476 iovdd.n475 0.00900667
R1575 iovdd.n551 iovdd.n550 0.00871333
R1576 iovdd.n462 iovdd.n461 0.00871333
R1577 iovdd.n562 iovdd.n224 0.00856667
R1578 iovdd.n667 iovdd 0.00851289
R1579 iovdd.n506 iovdd.n505 0.00827333
R1580 iovdd.n448 iovdd.n447 0.00798
R1581 iovdd.n647 iovdd.n646 0.00783333
R1582 iovdd.n646 iovdd.n645 0.00783333
R1583 iovdd.n666 iovdd.n82 0.00783333
R1584 iovdd.n662 iovdd.n82 0.00783333
R1585 iovdd.n545 iovdd.n544 0.00783333
R1586 iovdd.n469 iovdd.n468 0.00783333
R1587 iovdd.n544 iovdd.n543 0.00754
R1588 iovdd.n470 iovdd.n469 0.00754
R1589 iovdd.n701 iovdd.n700 0.00740196
R1590 iovdd.n702 iovdd.n701 0.00740196
R1591 iovdd.n702 iovdd.n681 0.00740196
R1592 iovdd.n715 iovdd.n681 0.00740196
R1593 iovdd.n716 iovdd.n715 0.00740196
R1594 iovdd.n717 iovdd.n716 0.00740196
R1595 iovdd.n718 iovdd.n717 0.00740196
R1596 iovdd.n728 iovdd.n718 0.00740196
R1597 iovdd.n729 iovdd.n728 0.00740196
R1598 iovdd.n730 iovdd.n729 0.00740196
R1599 iovdd.n731 iovdd.n730 0.00740196
R1600 iovdd.n741 iovdd.n731 0.00740196
R1601 iovdd.n742 iovdd.n741 0.00740196
R1602 iovdd.n743 iovdd.n742 0.00740196
R1603 iovdd.n744 iovdd.n743 0.00740196
R1604 iovdd.n749 iovdd.n744 0.00740196
R1605 iovdd.n807 iovdd.n749 0.00740196
R1606 iovdd.n808 iovdd.n807 0.00740196
R1607 iovdd.n819 iovdd.n808 0.00740196
R1608 iovdd.n820 iovdd.n819 0.00740196
R1609 iovdd.n821 iovdd.n820 0.00740196
R1610 iovdd.n822 iovdd.n821 0.00740196
R1611 iovdd.n832 iovdd.n822 0.00740196
R1612 iovdd.n833 iovdd.n832 0.00740196
R1613 iovdd.n834 iovdd.n833 0.00740196
R1614 iovdd.n835 iovdd.n834 0.00740196
R1615 iovdd.n844 iovdd.n835 0.00740196
R1616 iovdd.n845 iovdd.n844 0.00740196
R1617 iovdd.n846 iovdd.n845 0.00740196
R1618 iovdd.n847 iovdd.n846 0.00740196
R1619 iovdd.n858 iovdd.n847 0.00740196
R1620 iovdd.n859 iovdd.n858 0.00740196
R1621 iovdd.n860 iovdd.n859 0.00740196
R1622 iovdd.n861 iovdd.n860 0.00740196
R1623 iovdd.n864 iovdd.n861 0.00740196
R1624 iovdd.n865 iovdd.n864 0.00740196
R1625 iovdd.n865 iovdd 0.00740196
R1626 iovdd.n699 iovdd.n691 0.00740196
R1627 iovdd.n699 iovdd.n689 0.00740196
R1628 iovdd.n703 iovdd.n689 0.00740196
R1629 iovdd.n703 iovdd.n682 0.00740196
R1630 iovdd.n714 iovdd.n682 0.00740196
R1631 iovdd.n714 iovdd.n680 0.00740196
R1632 iovdd.n951 iovdd.n680 0.00740196
R1633 iovdd.n951 iovdd.n950 0.00740196
R1634 iovdd.n950 iovdd.n719 0.00740196
R1635 iovdd.n727 iovdd.n719 0.00740196
R1636 iovdd.n940 iovdd.n727 0.00740196
R1637 iovdd.n940 iovdd.n939 0.00740196
R1638 iovdd.n939 iovdd.n732 0.00740196
R1639 iovdd.n740 iovdd.n732 0.00740196
R1640 iovdd.n929 iovdd.n740 0.00740196
R1641 iovdd.n929 iovdd.n928 0.00740196
R1642 iovdd.n928 iovdd.n745 0.00740196
R1643 iovdd.n919 iovdd.n745 0.00740196
R1644 iovdd.n919 iovdd.n918 0.00740196
R1645 iovdd.n918 iovdd.n809 0.00740196
R1646 iovdd.n818 iovdd.n809 0.00740196
R1647 iovdd.n908 iovdd.n818 0.00740196
R1648 iovdd.n908 iovdd.n907 0.00740196
R1649 iovdd.n907 iovdd.n823 0.00740196
R1650 iovdd.n831 iovdd.n823 0.00740196
R1651 iovdd.n897 iovdd.n831 0.00740196
R1652 iovdd.n897 iovdd.n896 0.00740196
R1653 iovdd.n896 iovdd.n836 0.00740196
R1654 iovdd.n843 iovdd.n836 0.00740196
R1655 iovdd.n886 iovdd.n843 0.00740196
R1656 iovdd.n886 iovdd.n885 0.00740196
R1657 iovdd.n885 iovdd.n848 0.00740196
R1658 iovdd.n857 iovdd.n848 0.00740196
R1659 iovdd.n875 iovdd.n857 0.00740196
R1660 iovdd.n875 iovdd.n874 0.00740196
R1661 iovdd.n874 iovdd.n862 0.00740196
R1662 iovdd.n866 iovdd.n862 0.00740196
R1663 iovdd.n971 iovdd.n962 0.00740196
R1664 iovdd.n984 iovdd.n962 0.00740196
R1665 iovdd.n985 iovdd.n984 0.00740196
R1666 iovdd.n986 iovdd.n985 0.00740196
R1667 iovdd.n986 iovdd.n71 0.00740196
R1668 iovdd.n1000 iovdd.n71 0.00740196
R1669 iovdd.n1001 iovdd.n1000 0.00740196
R1670 iovdd.n1002 iovdd.n1001 0.00740196
R1671 iovdd.n1002 iovdd.n62 0.00740196
R1672 iovdd.n1015 iovdd.n62 0.00740196
R1673 iovdd.n1016 iovdd.n1015 0.00740196
R1674 iovdd.n1017 iovdd.n1016 0.00740196
R1675 iovdd.n1017 iovdd.n53 0.00740196
R1676 iovdd.n1030 iovdd.n53 0.00740196
R1677 iovdd.n1031 iovdd.n1030 0.00740196
R1678 iovdd.n1032 iovdd.n1031 0.00740196
R1679 iovdd.n1032 iovdd.n42 0.00740196
R1680 iovdd.n1046 iovdd.n42 0.00740196
R1681 iovdd.n1047 iovdd.n1046 0.00740196
R1682 iovdd.n1048 iovdd.n1047 0.00740196
R1683 iovdd.n1048 iovdd.n33 0.00740196
R1684 iovdd.n1061 iovdd.n33 0.00740196
R1685 iovdd.n1062 iovdd.n1061 0.00740196
R1686 iovdd.n1063 iovdd.n1062 0.00740196
R1687 iovdd.n1063 iovdd.n24 0.00740196
R1688 iovdd.n1076 iovdd.n24 0.00740196
R1689 iovdd.n1077 iovdd.n1076 0.00740196
R1690 iovdd.n1078 iovdd.n1077 0.00740196
R1691 iovdd.n1078 iovdd.n13 0.00740196
R1692 iovdd.n1092 iovdd.n13 0.00740196
R1693 iovdd.n1093 iovdd.n1092 0.00740196
R1694 iovdd.n1094 iovdd.n1093 0.00740196
R1695 iovdd.n1094 iovdd.n4 0.00740196
R1696 iovdd.n1107 iovdd.n4 0.00740196
R1697 iovdd.n972 iovdd.n969 0.00740196
R1698 iovdd.n972 iovdd.n963 0.00740196
R1699 iovdd.n983 iovdd.n963 0.00740196
R1700 iovdd.n983 iovdd.n961 0.00740196
R1701 iovdd.n987 iovdd.n961 0.00740196
R1702 iovdd.n987 iovdd.n72 0.00740196
R1703 iovdd.n999 iovdd.n72 0.00740196
R1704 iovdd.n999 iovdd.n70 0.00740196
R1705 iovdd.n1003 iovdd.n70 0.00740196
R1706 iovdd.n1003 iovdd.n63 0.00740196
R1707 iovdd.n1014 iovdd.n63 0.00740196
R1708 iovdd.n1014 iovdd.n61 0.00740196
R1709 iovdd.n1018 iovdd.n61 0.00740196
R1710 iovdd.n1018 iovdd.n54 0.00740196
R1711 iovdd.n1029 iovdd.n54 0.00740196
R1712 iovdd.n1029 iovdd.n52 0.00740196
R1713 iovdd.n1033 iovdd.n52 0.00740196
R1714 iovdd.n1033 iovdd.n43 0.00740196
R1715 iovdd.n1045 iovdd.n43 0.00740196
R1716 iovdd.n1045 iovdd.n41 0.00740196
R1717 iovdd.n1049 iovdd.n41 0.00740196
R1718 iovdd.n1049 iovdd.n34 0.00740196
R1719 iovdd.n1060 iovdd.n34 0.00740196
R1720 iovdd.n1060 iovdd.n32 0.00740196
R1721 iovdd.n1064 iovdd.n32 0.00740196
R1722 iovdd.n1064 iovdd.n25 0.00740196
R1723 iovdd.n1075 iovdd.n25 0.00740196
R1724 iovdd.n1075 iovdd.n23 0.00740196
R1725 iovdd.n1079 iovdd.n23 0.00740196
R1726 iovdd.n1079 iovdd.n14 0.00740196
R1727 iovdd.n1091 iovdd.n14 0.00740196
R1728 iovdd.n1091 iovdd.n12 0.00740196
R1729 iovdd.n1095 iovdd.n12 0.00740196
R1730 iovdd.n1095 iovdd.n5 0.00740196
R1731 iovdd.n1106 iovdd.n5 0.00740196
R1732 iovdd.n1106 iovdd.n3 0.00740196
R1733 iovdd.n447 iovdd.n446 0.00739333
R1734 iovdd.n505 iovdd.n504 0.0071
R1735 iovdd.n659 iovdd.n658 0.00696745
R1736 iovdd.n656 iovdd.n655 0.00696745
R1737 iovdd.n653 iovdd.n652 0.00696745
R1738 iovdd.n650 iovdd.n649 0.00696745
R1739 iovdd.n643 iovdd.n642 0.00696745
R1740 iovdd.n640 iovdd.n639 0.00696745
R1741 iovdd.n637 iovdd.n636 0.00696745
R1742 iovdd.n634 iovdd.n633 0.00696745
R1743 iovdd.n660 iovdd.n659 0.00696745
R1744 iovdd.n657 iovdd.n656 0.00696745
R1745 iovdd.n654 iovdd.n653 0.00696745
R1746 iovdd.n651 iovdd.n650 0.00696745
R1747 iovdd.n642 iovdd.n641 0.00696745
R1748 iovdd.n639 iovdd.n638 0.00696745
R1749 iovdd.n636 iovdd.n635 0.00696745
R1750 iovdd.n633 iovdd.n632 0.00696745
R1751 iovdd.n559 iovdd.n224 0.00680667
R1752 iovdd.n551 iovdd.n232 0.00666
R1753 iovdd.n461 iovdd.n348 0.00666
R1754 iovdd.n536 iovdd.n253 0.00636667
R1755 iovdd.n476 iovdd.n327 0.00636667
R1756 iovdd.n572 iovdd.n215 0.00622
R1757 iovdd.n626 iovdd.n108 0.00607333
R1758 iovdd.n804 iovdd.n750 0.00603377
R1759 iovdd.n629 iovdd.n18 0.006
R1760 iovdd.n292 iovdd.n291 0.00592667
R1761 iovdd.n363 iovdd.n362 0.00563333
R1762 iovdd.n556 iovdd.n555 0.00548667
R1763 iovdd.n458 iovdd.n457 0.00548667
R1764 iovdd.n533 iovdd.n532 0.00519333
R1765 iovdd.n480 iovdd.n479 0.00519333
R1766 iovdd.n438 iovdd.n387 0.00504667
R1767 iovdd.n596 iovdd.n142 0.0049
R1768 iovdd.n617 iovdd.n111 0.0049
R1769 iovdd.n494 iovdd.n493 0.00475333
R1770 iovdd.n244 iovdd.n243 0.00446
R1771 iovdd.n691 iovdd.n690 0.00442211
R1772 iovdd.n1108 iovdd.n3 0.00442211
R1773 iovdd.n970 iovdd.n969 0.00442211
R1774 iovdd.n225 iovdd.n218 0.00431333
R1775 iovdd.n451 iovdd.n450 0.00431333
R1776 iovdd.n629 iovdd 0.00416667
R1777 iovdd.n599 iovdd.n598 0.00416667
R1778 iovdd.n526 iovdd.n525 0.00402
R1779 iovdd.n318 iovdd.n311 0.00402
R1780 iovdd.n693 iovdd.n692 0.00395098
R1781 iovdd.n696 iovdd.n692 0.00395098
R1782 iovdd.n698 iovdd.n696 0.00395098
R1783 iovdd.n698 iovdd.n697 0.00395098
R1784 iovdd.n697 iovdd.n687 0.00395098
R1785 iovdd.n705 iovdd.n687 0.00395098
R1786 iovdd.n705 iovdd.n704 0.00395098
R1787 iovdd.n704 iovdd.n688 0.00395098
R1788 iovdd.n688 iovdd.n683 0.00395098
R1789 iovdd.n711 iovdd.n683 0.00395098
R1790 iovdd.n713 iovdd.n711 0.00395098
R1791 iovdd.n713 iovdd.n712 0.00395098
R1792 iovdd.n712 iovdd.n678 0.00395098
R1793 iovdd.n953 iovdd.n678 0.00395098
R1794 iovdd.n953 iovdd.n952 0.00395098
R1795 iovdd.n952 iovdd.n679 0.00395098
R1796 iovdd.n949 iovdd.n679 0.00395098
R1797 iovdd.n949 iovdd.n948 0.00395098
R1798 iovdd.n948 iovdd.n720 0.00395098
R1799 iovdd.n724 iovdd.n720 0.00395098
R1800 iovdd.n725 iovdd.n724 0.00395098
R1801 iovdd.n942 iovdd.n725 0.00395098
R1802 iovdd.n942 iovdd.n941 0.00395098
R1803 iovdd.n941 iovdd.n726 0.00395098
R1804 iovdd.n938 iovdd.n726 0.00395098
R1805 iovdd.n938 iovdd.n937 0.00395098
R1806 iovdd.n937 iovdd.n733 0.00395098
R1807 iovdd.n737 iovdd.n733 0.00395098
R1808 iovdd.n738 iovdd.n737 0.00395098
R1809 iovdd.n931 iovdd.n738 0.00395098
R1810 iovdd.n931 iovdd.n930 0.00395098
R1811 iovdd.n930 iovdd.n739 0.00395098
R1812 iovdd.n927 iovdd.n739 0.00395098
R1813 iovdd.n927 iovdd.n926 0.00395098
R1814 iovdd.n926 iovdd.n746 0.00395098
R1815 iovdd.n921 iovdd.n746 0.00395098
R1816 iovdd.n921 iovdd.n920 0.00395098
R1817 iovdd.n920 iovdd.n748 0.00395098
R1818 iovdd.n917 iovdd.n748 0.00395098
R1819 iovdd.n917 iovdd.n916 0.00395098
R1820 iovdd.n916 iovdd.n810 0.00395098
R1821 iovdd.n815 iovdd.n810 0.00395098
R1822 iovdd.n816 iovdd.n815 0.00395098
R1823 iovdd.n910 iovdd.n816 0.00395098
R1824 iovdd.n910 iovdd.n909 0.00395098
R1825 iovdd.n909 iovdd.n817 0.00395098
R1826 iovdd.n906 iovdd.n817 0.00395098
R1827 iovdd.n906 iovdd.n905 0.00395098
R1828 iovdd.n905 iovdd.n824 0.00395098
R1829 iovdd.n828 iovdd.n824 0.00395098
R1830 iovdd.n829 iovdd.n828 0.00395098
R1831 iovdd.n899 iovdd.n829 0.00395098
R1832 iovdd.n899 iovdd.n898 0.00395098
R1833 iovdd.n898 iovdd.n830 0.00395098
R1834 iovdd.n895 iovdd.n830 0.00395098
R1835 iovdd.n895 iovdd.n894 0.00395098
R1836 iovdd.n894 iovdd.n837 0.00395098
R1837 iovdd.n840 iovdd.n837 0.00395098
R1838 iovdd.n841 iovdd.n840 0.00395098
R1839 iovdd.n888 iovdd.n841 0.00395098
R1840 iovdd.n888 iovdd.n887 0.00395098
R1841 iovdd.n887 iovdd.n842 0.00395098
R1842 iovdd.n884 iovdd.n842 0.00395098
R1843 iovdd.n884 iovdd.n883 0.00395098
R1844 iovdd.n883 iovdd.n849 0.00395098
R1845 iovdd.n854 iovdd.n849 0.00395098
R1846 iovdd.n855 iovdd.n854 0.00395098
R1847 iovdd.n877 iovdd.n855 0.00395098
R1848 iovdd.n877 iovdd.n876 0.00395098
R1849 iovdd.n876 iovdd.n856 0.00395098
R1850 iovdd.n873 iovdd.n856 0.00395098
R1851 iovdd.n873 iovdd.n872 0.00395098
R1852 iovdd.n872 iovdd.n863 0.00395098
R1853 iovdd.n867 iovdd.n863 0.00395098
R1854 iovdd.n967 iovdd.n966 0.00395098
R1855 iovdd.n974 iovdd.n967 0.00395098
R1856 iovdd.n974 iovdd.n973 0.00395098
R1857 iovdd.n973 iovdd.n968 0.00395098
R1858 iovdd.n968 iovdd.n964 0.00395098
R1859 iovdd.n980 iovdd.n964 0.00395098
R1860 iovdd.n982 iovdd.n980 0.00395098
R1861 iovdd.n982 iovdd.n981 0.00395098
R1862 iovdd.n981 iovdd.n959 0.00395098
R1863 iovdd.n989 iovdd.n959 0.00395098
R1864 iovdd.n989 iovdd.n988 0.00395098
R1865 iovdd.n988 iovdd.n960 0.00395098
R1866 iovdd.n960 iovdd.n73 0.00395098
R1867 iovdd.n996 iovdd.n73 0.00395098
R1868 iovdd.n998 iovdd.n996 0.00395098
R1869 iovdd.n998 iovdd.n997 0.00395098
R1870 iovdd.n997 iovdd.n68 0.00395098
R1871 iovdd.n1005 iovdd.n68 0.00395098
R1872 iovdd.n1005 iovdd.n1004 0.00395098
R1873 iovdd.n1004 iovdd.n69 0.00395098
R1874 iovdd.n69 iovdd.n64 0.00395098
R1875 iovdd.n1011 iovdd.n64 0.00395098
R1876 iovdd.n1013 iovdd.n1011 0.00395098
R1877 iovdd.n1013 iovdd.n1012 0.00395098
R1878 iovdd.n1012 iovdd.n59 0.00395098
R1879 iovdd.n1020 iovdd.n59 0.00395098
R1880 iovdd.n1020 iovdd.n1019 0.00395098
R1881 iovdd.n1019 iovdd.n60 0.00395098
R1882 iovdd.n60 iovdd.n55 0.00395098
R1883 iovdd.n1026 iovdd.n55 0.00395098
R1884 iovdd.n1028 iovdd.n1026 0.00395098
R1885 iovdd.n1028 iovdd.n1027 0.00395098
R1886 iovdd.n1027 iovdd.n50 0.00395098
R1887 iovdd.n1035 iovdd.n50 0.00395098
R1888 iovdd.n1035 iovdd.n1034 0.00395098
R1889 iovdd.n1034 iovdd.n51 0.00395098
R1890 iovdd.n51 iovdd.n44 0.00395098
R1891 iovdd.n1042 iovdd.n44 0.00395098
R1892 iovdd.n1044 iovdd.n1042 0.00395098
R1893 iovdd.n1044 iovdd.n1043 0.00395098
R1894 iovdd.n1043 iovdd.n39 0.00395098
R1895 iovdd.n1051 iovdd.n39 0.00395098
R1896 iovdd.n1051 iovdd.n1050 0.00395098
R1897 iovdd.n1050 iovdd.n40 0.00395098
R1898 iovdd.n40 iovdd.n35 0.00395098
R1899 iovdd.n1057 iovdd.n35 0.00395098
R1900 iovdd.n1059 iovdd.n1057 0.00395098
R1901 iovdd.n1059 iovdd.n1058 0.00395098
R1902 iovdd.n1058 iovdd.n30 0.00395098
R1903 iovdd.n1066 iovdd.n30 0.00395098
R1904 iovdd.n1066 iovdd.n1065 0.00395098
R1905 iovdd.n1065 iovdd.n31 0.00395098
R1906 iovdd.n31 iovdd.n26 0.00395098
R1907 iovdd.n1072 iovdd.n26 0.00395098
R1908 iovdd.n1074 iovdd.n1072 0.00395098
R1909 iovdd.n1074 iovdd.n1073 0.00395098
R1910 iovdd.n1073 iovdd.n21 0.00395098
R1911 iovdd.n1081 iovdd.n21 0.00395098
R1912 iovdd.n1081 iovdd.n1080 0.00395098
R1913 iovdd.n1080 iovdd.n22 0.00395098
R1914 iovdd.n22 iovdd.n15 0.00395098
R1915 iovdd.n1088 iovdd.n15 0.00395098
R1916 iovdd.n1090 iovdd.n1088 0.00395098
R1917 iovdd.n1090 iovdd.n1089 0.00395098
R1918 iovdd.n1089 iovdd.n10 0.00395098
R1919 iovdd.n1097 iovdd.n10 0.00395098
R1920 iovdd.n1097 iovdd.n1096 0.00395098
R1921 iovdd.n1096 iovdd.n11 0.00395098
R1922 iovdd.n11 iovdd.n6 0.00395098
R1923 iovdd.n1103 iovdd.n6 0.00395098
R1924 iovdd.n1105 iovdd.n1103 0.00395098
R1925 iovdd.n1105 iovdd.n1104 0.00395098
R1926 iovdd.n1104 iovdd.n2 0.00395098
R1927 iovdd.n1109 iovdd.n2 0.00395098
R1928 iovdd.n582 iovdd.n581 0.00387333
R1929 iovdd.n606 iovdd.n137 0.00383939
R1930 iovdd.n176 iovdd.n166 0.00372667
R1931 iovdd.n410 iovdd.n409 0.00372667
R1932 iovdd.n662 iovdd.n46 0.00358
R1933 iovdd.n523 iovdd.n522 0.00358
R1934 iovdd.n647 iovdd.n46 0.00354333
R1935 iovdd.n1039 iovdd.n47 0.00350055
R1936 iovdd.n993 iovdd.n956 0.00350055
R1937 iovdd.n1085 iovdd.n17 0.00350055
R1938 iovdd.n466 iovdd.n465 0.00328667
R1939 iovdd.n570 iovdd.n216 0.00314
R1940 iovdd.n443 iovdd.n372 0.00314
R1941 iovdd.n614 iovdd.n613 0.00299333
R1942 iovdd.n518 iovdd.n277 0.00284667
R1943 iovdd.n310 iovdd.n303 0.00284667
R1944 iovdd.n429 iovdd.n428 0.0027
R1945 iovdd.n1110 iovdd 0.00261765
R1946 iovdd.n185 iovdd.n164 0.00255333
R1947 iovdd.n405 iovdd.n398 0.00255333
R1948 iovdd.n483 iovdd.n317 0.00240667
R1949 iovdd.n541 iovdd.n540 0.00211333
R1950 iovdd.n577 iovdd.n576 0.00196667
R1951 iovdd.n440 iovdd.n439 0.00196667
R1952 iovdd.n869 iovdd 0.00196667
R1953 iovdd iovdd.n1111 0.00196667
R1954 iovdd.n695 iovdd.n686 0.00191176
R1955 iovdd.n706 iovdd.n686 0.00191176
R1956 iovdd.n706 iovdd.n684 0.00191176
R1957 iovdd.n710 iovdd.n684 0.00191176
R1958 iovdd.n710 iovdd.n676 0.00191176
R1959 iovdd.n954 iovdd.n676 0.00191176
R1960 iovdd.n954 iovdd.n677 0.00191176
R1961 iovdd.n947 iovdd.n677 0.00191176
R1962 iovdd.n947 iovdd.n721 0.00191176
R1963 iovdd.n943 iovdd.n721 0.00191176
R1964 iovdd.n943 iovdd.n723 0.00191176
R1965 iovdd.n936 iovdd.n723 0.00191176
R1966 iovdd.n936 iovdd.n734 0.00191176
R1967 iovdd.n932 iovdd.n734 0.00191176
R1968 iovdd.n932 iovdd.n736 0.00191176
R1969 iovdd.n925 iovdd.n736 0.00191176
R1970 iovdd.n925 iovdd.n922 0.00191176
R1971 iovdd.n922 iovdd.n747 0.00191176
R1972 iovdd.n915 iovdd.n747 0.00191176
R1973 iovdd.n915 iovdd.n811 0.00191176
R1974 iovdd.n911 iovdd.n811 0.00191176
R1975 iovdd.n911 iovdd.n814 0.00191176
R1976 iovdd.n904 iovdd.n814 0.00191176
R1977 iovdd.n904 iovdd.n825 0.00191176
R1978 iovdd.n900 iovdd.n825 0.00191176
R1979 iovdd.n900 iovdd.n827 0.00191176
R1980 iovdd.n893 iovdd.n827 0.00191176
R1981 iovdd.n893 iovdd.n838 0.00191176
R1982 iovdd.n889 iovdd.n838 0.00191176
R1983 iovdd.n889 iovdd.n839 0.00191176
R1984 iovdd.n882 iovdd.n839 0.00191176
R1985 iovdd.n882 iovdd.n850 0.00191176
R1986 iovdd.n878 iovdd.n850 0.00191176
R1987 iovdd.n878 iovdd.n853 0.00191176
R1988 iovdd.n871 iovdd.n853 0.00191176
R1989 iovdd.n871 iovdd.n868 0.00191176
R1990 iovdd.n975 iovdd.n965 0.00191176
R1991 iovdd.n979 iovdd.n965 0.00191176
R1992 iovdd.n979 iovdd.n958 0.00191176
R1993 iovdd.n990 iovdd.n958 0.00191176
R1994 iovdd.n990 iovdd.n74 0.00191176
R1995 iovdd.n995 iovdd.n74 0.00191176
R1996 iovdd.n995 iovdd.n67 0.00191176
R1997 iovdd.n1006 iovdd.n67 0.00191176
R1998 iovdd.n1006 iovdd.n65 0.00191176
R1999 iovdd.n1010 iovdd.n65 0.00191176
R2000 iovdd.n1010 iovdd.n58 0.00191176
R2001 iovdd.n1021 iovdd.n58 0.00191176
R2002 iovdd.n1021 iovdd.n56 0.00191176
R2003 iovdd.n1025 iovdd.n56 0.00191176
R2004 iovdd.n1025 iovdd.n49 0.00191176
R2005 iovdd.n1036 iovdd.n49 0.00191176
R2006 iovdd.n1036 iovdd.n45 0.00191176
R2007 iovdd.n1041 iovdd.n45 0.00191176
R2008 iovdd.n1041 iovdd.n38 0.00191176
R2009 iovdd.n1052 iovdd.n38 0.00191176
R2010 iovdd.n1052 iovdd.n36 0.00191176
R2011 iovdd.n1056 iovdd.n36 0.00191176
R2012 iovdd.n1056 iovdd.n29 0.00191176
R2013 iovdd.n1067 iovdd.n29 0.00191176
R2014 iovdd.n1067 iovdd.n27 0.00191176
R2015 iovdd.n1071 iovdd.n27 0.00191176
R2016 iovdd.n1071 iovdd.n20 0.00191176
R2017 iovdd.n1082 iovdd.n20 0.00191176
R2018 iovdd.n1082 iovdd.n16 0.00191176
R2019 iovdd.n1087 iovdd.n16 0.00191176
R2020 iovdd.n1087 iovdd.n9 0.00191176
R2021 iovdd.n1098 iovdd.n9 0.00191176
R2022 iovdd.n1098 iovdd.n7 0.00191176
R2023 iovdd.n1102 iovdd.n7 0.00191176
R2024 iovdd.n1102 iovdd.n1 0.00191176
R2025 iovdd.n1110 iovdd.n1 0.00191176
R2026 iovdd.n181 iovdd.n180 0.00182
R2027 iovdd.n695 iovdd.n694 0.0016983
R2028 iovdd.n976 iovdd.n975 0.0016983
R2029 iovdd.n515 iovdd.n514 0.00167333
R2030 iovdd.n501 iovdd.n301 0.00167333
R2031 iovdd.n195 iovdd.n194 0.00152667
R2032 iovdd.n707 iovdd.n685 0.00147778
R2033 iovdd.n708 iovdd.n707 0.00147778
R2034 iovdd.n709 iovdd.n708 0.00147778
R2035 iovdd.n709 iovdd.n674 0.00147778
R2036 iovdd.n955 iovdd.n675 0.00147778
R2037 iovdd.n946 iovdd.n675 0.00147778
R2038 iovdd.n946 iovdd.n945 0.00147778
R2039 iovdd.n945 iovdd.n944 0.00147778
R2040 iovdd.n944 iovdd.n722 0.00147778
R2041 iovdd.n935 iovdd.n722 0.00147778
R2042 iovdd.n935 iovdd.n934 0.00147778
R2043 iovdd.n934 iovdd.n933 0.00147778
R2044 iovdd.n933 iovdd.n735 0.00147778
R2045 iovdd.n924 iovdd.n735 0.00147778
R2046 iovdd.n924 iovdd.n923 0.00147778
R2047 iovdd.n914 iovdd.n812 0.00147778
R2048 iovdd.n914 iovdd.n913 0.00147778
R2049 iovdd.n913 iovdd.n912 0.00147778
R2050 iovdd.n912 iovdd.n813 0.00147778
R2051 iovdd.n903 iovdd.n813 0.00147778
R2052 iovdd.n903 iovdd.n902 0.00147778
R2053 iovdd.n902 iovdd.n901 0.00147778
R2054 iovdd.n901 iovdd.n826 0.00147778
R2055 iovdd.n892 iovdd.n826 0.00147778
R2056 iovdd.n892 iovdd.n891 0.00147778
R2057 iovdd.n891 iovdd.n890 0.00147778
R2058 iovdd.n881 iovdd.n851 0.00147778
R2059 iovdd.n881 iovdd.n880 0.00147778
R2060 iovdd.n880 iovdd.n879 0.00147778
R2061 iovdd.n879 iovdd.n852 0.00147778
R2062 iovdd.n870 iovdd.n852 0.00147778
R2063 iovdd.n870 iovdd.n869 0.00147778
R2064 iovdd.n978 iovdd.n977 0.00147778
R2065 iovdd.n978 iovdd.n957 0.00147778
R2066 iovdd.n991 iovdd.n957 0.00147778
R2067 iovdd.n992 iovdd.n991 0.00147778
R2068 iovdd.n994 iovdd.n66 0.00147778
R2069 iovdd.n1007 iovdd.n66 0.00147778
R2070 iovdd.n1008 iovdd.n1007 0.00147778
R2071 iovdd.n1009 iovdd.n1008 0.00147778
R2072 iovdd.n1009 iovdd.n57 0.00147778
R2073 iovdd.n1022 iovdd.n57 0.00147778
R2074 iovdd.n1023 iovdd.n1022 0.00147778
R2075 iovdd.n1024 iovdd.n1023 0.00147778
R2076 iovdd.n1024 iovdd.n48 0.00147778
R2077 iovdd.n1037 iovdd.n48 0.00147778
R2078 iovdd.n1038 iovdd.n1037 0.00147778
R2079 iovdd.n1040 iovdd.n37 0.00147778
R2080 iovdd.n1053 iovdd.n37 0.00147778
R2081 iovdd.n1054 iovdd.n1053 0.00147778
R2082 iovdd.n1055 iovdd.n1054 0.00147778
R2083 iovdd.n1055 iovdd.n28 0.00147778
R2084 iovdd.n1068 iovdd.n28 0.00147778
R2085 iovdd.n1069 iovdd.n1068 0.00147778
R2086 iovdd.n1070 iovdd.n1069 0.00147778
R2087 iovdd.n1070 iovdd.n19 0.00147778
R2088 iovdd.n1083 iovdd.n19 0.00147778
R2089 iovdd.n1084 iovdd.n1083 0.00147778
R2090 iovdd.n1086 iovdd.n8 0.00147778
R2091 iovdd.n1099 iovdd.n8 0.00147778
R2092 iovdd.n1100 iovdd.n1099 0.00147778
R2093 iovdd.n1101 iovdd.n1100 0.00147778
R2094 iovdd.n1101 iovdd.n0 0.00147778
R2095 iovdd.n1111 iovdd.n0 0.00147778
R2096 iovdd.n46 iovdd 0.00140016
R2097 iovdd.n18 iovdd 0.00140016
R2098 iovdd.n192 iovdd.n157 0.00138
R2099 iovdd.n425 iovdd.n396 0.00138
R2100 iovdd.n956 iovdd.n674 0.001314
R2101 iovdd.n851 iovdd.n17 0.001314
R2102 iovdd.n993 iovdd.n992 0.001314
R2103 iovdd.n1086 iovdd.n1085 0.001314
R2104 iovdd.n268 iovdd.n267 0.00123333
R2105 iovdd.n645 iovdd.n18 0.00112333
R2106 iovdd.n667 iovdd.n666 0.00112333
R2107 iovdd.n606 iovdd.n138 0.00100123
R2108 iovdd.n923 iovdd.n47 0.000991333
R2109 iovdd.n1039 iovdd.n1038 0.000991333
R2110 iovdd.n812 iovdd.n47 0.000986444
R2111 iovdd.n1040 iovdd.n1039 0.000986444
R2112 iovdd.n339 iovdd.n338 0.00094
R2113 iovdd.n592 iovdd.n591 0.000825926
R2114 iovdd.n591 iovdd.n590 0.000825926
R2115 iovdd.n590 iovdd.n150 0.000825926
R2116 iovdd.n150 iovdd.n75 0.000825926
R2117 iovdd.n673 iovdd.n76 0.000825926
R2118 iovdd.n669 iovdd.n76 0.000825926
R2119 iovdd.n669 iovdd.n668 0.000825926
R2120 iovdd.n668 iovdd.n667 0.000798222
R2121 iovdd.n584 iovdd.n154 0.000793333
R2122 iovdd.n433 iovdd.n432 0.000793333
R2123 iovdd.n993 iovdd.n673 0.000717556
R2124 iovdd.n956 iovdd.n955 0.000663778
R2125 iovdd.n890 iovdd.n17 0.000663778
R2126 iovdd.n994 iovdd.n993 0.000663778
R2127 iovdd.n1085 iovdd.n1084 0.000663778
R2128 iovdd.n418 iovdd.n417 0.000646667
R2129 iovdd.n993 iovdd.n75 0.00060837
R2130 iovdd.n592 iovdd.n149 0.000581482
R2131 iovss.n87 iovss.n85 0.826084
R2132 iovss.n186 iovss.n1 0.826084
R2133 iovss.n86 iovss.n81 0.818682
R2134 iovss.n95 iovss.n80 0.818682
R2135 iovss.n96 iovss.n79 0.818682
R2136 iovss.n78 iovss.n74 0.818682
R2137 iovss.n103 iovss.n73 0.818682
R2138 iovss.n104 iovss.n72 0.818682
R2139 iovss.n71 iovss.n67 0.818682
R2140 iovss.n111 iovss.n66 0.818682
R2141 iovss.n112 iovss.n65 0.818682
R2142 iovss.n64 iovss.n60 0.818682
R2143 iovss.n119 iovss.n59 0.818682
R2144 iovss.n120 iovss.n58 0.818682
R2145 iovss.n57 iovss.n53 0.818682
R2146 iovss.n127 iovss.n52 0.818682
R2147 iovss.n128 iovss.n51 0.818682
R2148 iovss.n50 iovss.n46 0.818682
R2149 iovss.n135 iovss.n45 0.818682
R2150 iovss.n136 iovss.n44 0.818682
R2151 iovss.n43 iovss.n39 0.818682
R2152 iovss.n143 iovss.n38 0.818682
R2153 iovss.n144 iovss.n37 0.818682
R2154 iovss.n36 iovss.n32 0.818682
R2155 iovss.n151 iovss.n31 0.818682
R2156 iovss.n152 iovss.n30 0.818682
R2157 iovss.n29 iovss.n25 0.818682
R2158 iovss.n159 iovss.n24 0.818682
R2159 iovss.n160 iovss.n23 0.818682
R2160 iovss.n22 iovss.n18 0.818682
R2161 iovss.n167 iovss.n17 0.818682
R2162 iovss.n168 iovss.n16 0.818682
R2163 iovss.n15 iovss.n11 0.818682
R2164 iovss.n175 iovss.n10 0.818682
R2165 iovss.n176 iovss.n9 0.818682
R2166 iovss.n8 iovss.n4 0.818682
R2167 iovss.n183 iovss.n3 0.818682
R2168 iovss.n185 iovss.n184 0.818682
R2169 iovss.n183 iovss.n182 0.818682
R2170 iovss.n5 iovss.n4 0.818682
R2171 iovss.n177 iovss.n176 0.818682
R2172 iovss.n175 iovss.n174 0.818682
R2173 iovss.n12 iovss.n11 0.818682
R2174 iovss.n169 iovss.n168 0.818682
R2175 iovss.n167 iovss.n166 0.818682
R2176 iovss.n19 iovss.n18 0.818682
R2177 iovss.n161 iovss.n160 0.818682
R2178 iovss.n159 iovss.n158 0.818682
R2179 iovss.n26 iovss.n25 0.818682
R2180 iovss.n153 iovss.n152 0.818682
R2181 iovss.n151 iovss.n150 0.818682
R2182 iovss.n33 iovss.n32 0.818682
R2183 iovss.n145 iovss.n144 0.818682
R2184 iovss.n143 iovss.n142 0.818682
R2185 iovss.n40 iovss.n39 0.818682
R2186 iovss.n137 iovss.n136 0.818682
R2187 iovss.n135 iovss.n134 0.818682
R2188 iovss.n47 iovss.n46 0.818682
R2189 iovss.n129 iovss.n128 0.818682
R2190 iovss.n127 iovss.n126 0.818682
R2191 iovss.n54 iovss.n53 0.818682
R2192 iovss.n121 iovss.n120 0.818682
R2193 iovss.n119 iovss.n118 0.818682
R2194 iovss.n61 iovss.n60 0.818682
R2195 iovss.n113 iovss.n112 0.818682
R2196 iovss.n111 iovss.n110 0.818682
R2197 iovss.n68 iovss.n67 0.818682
R2198 iovss.n105 iovss.n104 0.818682
R2199 iovss.n103 iovss.n102 0.818682
R2200 iovss.n75 iovss.n74 0.818682
R2201 iovss.n97 iovss.n96 0.818682
R2202 iovss.n95 iovss.n94 0.818682
R2203 iovss.n82 iovss.n81 0.818682
R2204 iovss.n89 iovss.n88 0.818682
R2205 iovss.n3 iovss.n1 0.416993
R2206 iovss.n87 iovss.n86 0.416993
R2207 iovss.n85 iovss.n84 0.2005
R2208 iovss.n91 iovss.n90 0.2005
R2209 iovss.n93 iovss.n92 0.2005
R2210 iovss.n77 iovss.n76 0.2005
R2211 iovss.n99 iovss.n98 0.2005
R2212 iovss.n101 iovss.n100 0.2005
R2213 iovss.n70 iovss.n69 0.2005
R2214 iovss.n107 iovss.n106 0.2005
R2215 iovss.n109 iovss.n108 0.2005
R2216 iovss.n63 iovss.n62 0.2005
R2217 iovss.n115 iovss.n114 0.2005
R2218 iovss.n117 iovss.n116 0.2005
R2219 iovss.n56 iovss.n55 0.2005
R2220 iovss.n123 iovss.n122 0.2005
R2221 iovss.n125 iovss.n124 0.2005
R2222 iovss.n49 iovss.n48 0.2005
R2223 iovss.n131 iovss.n130 0.2005
R2224 iovss.n133 iovss.n132 0.2005
R2225 iovss.n42 iovss.n41 0.2005
R2226 iovss.n139 iovss.n138 0.2005
R2227 iovss.n141 iovss.n140 0.2005
R2228 iovss.n35 iovss.n34 0.2005
R2229 iovss.n147 iovss.n146 0.2005
R2230 iovss.n149 iovss.n148 0.2005
R2231 iovss.n28 iovss.n27 0.2005
R2232 iovss.n155 iovss.n154 0.2005
R2233 iovss.n157 iovss.n156 0.2005
R2234 iovss.n21 iovss.n20 0.2005
R2235 iovss.n163 iovss.n162 0.2005
R2236 iovss.n165 iovss.n164 0.2005
R2237 iovss.n14 iovss.n13 0.2005
R2238 iovss.n171 iovss.n170 0.2005
R2239 iovss.n173 iovss.n172 0.2005
R2240 iovss.n7 iovss.n6 0.2005
R2241 iovss.n179 iovss.n178 0.2005
R2242 iovss.n181 iovss.n180 0.2005
R2243 iovss.n2 iovss.n0 0.2005
R2244 iovss.n187 iovss.n186 0.2005
R2245 iovss iovss.n187 0.0778508
R2246 iovss.n83 iovss 0.0724109
R2247 iovss.n83 iovss 0.00862677
R2248 iovss.n84 iovss.n83 0.00808703
R2249 iovss.n8 iovss.n3 0.00740196
R2250 iovss.n9 iovss.n8 0.00740196
R2251 iovss.n10 iovss.n9 0.00740196
R2252 iovss.n15 iovss.n10 0.00740196
R2253 iovss.n16 iovss.n15 0.00740196
R2254 iovss.n17 iovss.n16 0.00740196
R2255 iovss.n22 iovss.n17 0.00740196
R2256 iovss.n23 iovss.n22 0.00740196
R2257 iovss.n24 iovss.n23 0.00740196
R2258 iovss.n29 iovss.n24 0.00740196
R2259 iovss.n30 iovss.n29 0.00740196
R2260 iovss.n31 iovss.n30 0.00740196
R2261 iovss.n36 iovss.n31 0.00740196
R2262 iovss.n37 iovss.n36 0.00740196
R2263 iovss.n38 iovss.n37 0.00740196
R2264 iovss.n43 iovss.n38 0.00740196
R2265 iovss.n44 iovss.n43 0.00740196
R2266 iovss.n45 iovss.n44 0.00740196
R2267 iovss.n50 iovss.n45 0.00740196
R2268 iovss.n51 iovss.n50 0.00740196
R2269 iovss.n52 iovss.n51 0.00740196
R2270 iovss.n57 iovss.n52 0.00740196
R2271 iovss.n58 iovss.n57 0.00740196
R2272 iovss.n59 iovss.n58 0.00740196
R2273 iovss.n64 iovss.n59 0.00740196
R2274 iovss.n65 iovss.n64 0.00740196
R2275 iovss.n66 iovss.n65 0.00740196
R2276 iovss.n71 iovss.n66 0.00740196
R2277 iovss.n72 iovss.n71 0.00740196
R2278 iovss.n73 iovss.n72 0.00740196
R2279 iovss.n78 iovss.n73 0.00740196
R2280 iovss.n79 iovss.n78 0.00740196
R2281 iovss.n80 iovss.n79 0.00740196
R2282 iovss.n86 iovss.n80 0.00740196
R2283 iovss.n184 iovss.n183 0.00740196
R2284 iovss.n183 iovss.n4 0.00740196
R2285 iovss.n176 iovss.n4 0.00740196
R2286 iovss.n176 iovss.n175 0.00740196
R2287 iovss.n175 iovss.n11 0.00740196
R2288 iovss.n168 iovss.n11 0.00740196
R2289 iovss.n168 iovss.n167 0.00740196
R2290 iovss.n167 iovss.n18 0.00740196
R2291 iovss.n160 iovss.n18 0.00740196
R2292 iovss.n160 iovss.n159 0.00740196
R2293 iovss.n159 iovss.n25 0.00740196
R2294 iovss.n152 iovss.n25 0.00740196
R2295 iovss.n152 iovss.n151 0.00740196
R2296 iovss.n151 iovss.n32 0.00740196
R2297 iovss.n144 iovss.n32 0.00740196
R2298 iovss.n144 iovss.n143 0.00740196
R2299 iovss.n143 iovss.n39 0.00740196
R2300 iovss.n136 iovss.n39 0.00740196
R2301 iovss.n136 iovss.n135 0.00740196
R2302 iovss.n135 iovss.n46 0.00740196
R2303 iovss.n128 iovss.n46 0.00740196
R2304 iovss.n128 iovss.n127 0.00740196
R2305 iovss.n127 iovss.n53 0.00740196
R2306 iovss.n120 iovss.n53 0.00740196
R2307 iovss.n120 iovss.n119 0.00740196
R2308 iovss.n119 iovss.n60 0.00740196
R2309 iovss.n112 iovss.n60 0.00740196
R2310 iovss.n112 iovss.n111 0.00740196
R2311 iovss.n111 iovss.n67 0.00740196
R2312 iovss.n104 iovss.n67 0.00740196
R2313 iovss.n104 iovss.n103 0.00740196
R2314 iovss.n103 iovss.n74 0.00740196
R2315 iovss.n96 iovss.n74 0.00740196
R2316 iovss.n96 iovss.n95 0.00740196
R2317 iovss.n95 iovss.n81 0.00740196
R2318 iovss.n88 iovss.n81 0.00740196
R2319 iovss.n88 iovss.n87 0.00442211
R2320 iovss.n184 iovss.n1 0.00442211
R2321 iovss.n186 iovss.n185 0.00395098
R2322 iovss.n185 iovss.n2 0.00395098
R2323 iovss.n182 iovss.n2 0.00395098
R2324 iovss.n182 iovss.n181 0.00395098
R2325 iovss.n181 iovss.n5 0.00395098
R2326 iovss.n178 iovss.n5 0.00395098
R2327 iovss.n178 iovss.n177 0.00395098
R2328 iovss.n177 iovss.n7 0.00395098
R2329 iovss.n174 iovss.n7 0.00395098
R2330 iovss.n174 iovss.n173 0.00395098
R2331 iovss.n173 iovss.n12 0.00395098
R2332 iovss.n170 iovss.n12 0.00395098
R2333 iovss.n170 iovss.n169 0.00395098
R2334 iovss.n169 iovss.n14 0.00395098
R2335 iovss.n166 iovss.n14 0.00395098
R2336 iovss.n166 iovss.n165 0.00395098
R2337 iovss.n165 iovss.n19 0.00395098
R2338 iovss.n162 iovss.n19 0.00395098
R2339 iovss.n162 iovss.n161 0.00395098
R2340 iovss.n161 iovss.n21 0.00395098
R2341 iovss.n158 iovss.n21 0.00395098
R2342 iovss.n158 iovss.n157 0.00395098
R2343 iovss.n157 iovss.n26 0.00395098
R2344 iovss.n154 iovss.n26 0.00395098
R2345 iovss.n154 iovss.n153 0.00395098
R2346 iovss.n153 iovss.n28 0.00395098
R2347 iovss.n150 iovss.n28 0.00395098
R2348 iovss.n150 iovss.n149 0.00395098
R2349 iovss.n149 iovss.n33 0.00395098
R2350 iovss.n146 iovss.n33 0.00395098
R2351 iovss.n146 iovss.n145 0.00395098
R2352 iovss.n145 iovss.n35 0.00395098
R2353 iovss.n142 iovss.n35 0.00395098
R2354 iovss.n142 iovss.n141 0.00395098
R2355 iovss.n141 iovss.n40 0.00395098
R2356 iovss.n138 iovss.n40 0.00395098
R2357 iovss.n138 iovss.n137 0.00395098
R2358 iovss.n137 iovss.n42 0.00395098
R2359 iovss.n134 iovss.n42 0.00395098
R2360 iovss.n134 iovss.n133 0.00395098
R2361 iovss.n133 iovss.n47 0.00395098
R2362 iovss.n130 iovss.n47 0.00395098
R2363 iovss.n130 iovss.n129 0.00395098
R2364 iovss.n129 iovss.n49 0.00395098
R2365 iovss.n126 iovss.n49 0.00395098
R2366 iovss.n126 iovss.n125 0.00395098
R2367 iovss.n125 iovss.n54 0.00395098
R2368 iovss.n122 iovss.n54 0.00395098
R2369 iovss.n122 iovss.n121 0.00395098
R2370 iovss.n121 iovss.n56 0.00395098
R2371 iovss.n118 iovss.n56 0.00395098
R2372 iovss.n118 iovss.n117 0.00395098
R2373 iovss.n117 iovss.n61 0.00395098
R2374 iovss.n114 iovss.n61 0.00395098
R2375 iovss.n114 iovss.n113 0.00395098
R2376 iovss.n113 iovss.n63 0.00395098
R2377 iovss.n110 iovss.n63 0.00395098
R2378 iovss.n110 iovss.n109 0.00395098
R2379 iovss.n109 iovss.n68 0.00395098
R2380 iovss.n106 iovss.n68 0.00395098
R2381 iovss.n106 iovss.n105 0.00395098
R2382 iovss.n105 iovss.n70 0.00395098
R2383 iovss.n102 iovss.n70 0.00395098
R2384 iovss.n102 iovss.n101 0.00395098
R2385 iovss.n101 iovss.n75 0.00395098
R2386 iovss.n98 iovss.n75 0.00395098
R2387 iovss.n98 iovss.n97 0.00395098
R2388 iovss.n97 iovss.n77 0.00395098
R2389 iovss.n94 iovss.n77 0.00395098
R2390 iovss.n94 iovss.n93 0.00395098
R2391 iovss.n93 iovss.n82 0.00395098
R2392 iovss.n90 iovss.n82 0.00395098
R2393 iovss.n90 iovss.n89 0.00395098
R2394 iovss.n89 iovss.n85 0.00395098
R2395 iovss.n187 iovss.n0 0.00191176
R2396 iovss.n180 iovss.n0 0.00191176
R2397 iovss.n180 iovss.n179 0.00191176
R2398 iovss.n179 iovss.n6 0.00191176
R2399 iovss.n172 iovss.n6 0.00191176
R2400 iovss.n172 iovss.n171 0.00191176
R2401 iovss.n171 iovss.n13 0.00191176
R2402 iovss.n164 iovss.n13 0.00191176
R2403 iovss.n164 iovss.n163 0.00191176
R2404 iovss.n163 iovss.n20 0.00191176
R2405 iovss.n156 iovss.n20 0.00191176
R2406 iovss.n156 iovss.n155 0.00191176
R2407 iovss.n155 iovss.n27 0.00191176
R2408 iovss.n148 iovss.n27 0.00191176
R2409 iovss.n148 iovss.n147 0.00191176
R2410 iovss.n147 iovss.n34 0.00191176
R2411 iovss.n140 iovss.n34 0.00191176
R2412 iovss.n140 iovss.n139 0.00191176
R2413 iovss.n139 iovss.n41 0.00191176
R2414 iovss.n132 iovss.n41 0.00191176
R2415 iovss.n132 iovss.n131 0.00191176
R2416 iovss.n131 iovss.n48 0.00191176
R2417 iovss.n124 iovss.n48 0.00191176
R2418 iovss.n124 iovss.n123 0.00191176
R2419 iovss.n123 iovss.n55 0.00191176
R2420 iovss.n116 iovss.n55 0.00191176
R2421 iovss.n116 iovss.n115 0.00191176
R2422 iovss.n115 iovss.n62 0.00191176
R2423 iovss.n108 iovss.n62 0.00191176
R2424 iovss.n108 iovss.n107 0.00191176
R2425 iovss.n107 iovss.n69 0.00191176
R2426 iovss.n100 iovss.n69 0.00191176
R2427 iovss.n100 iovss.n99 0.00191176
R2428 iovss.n99 iovss.n76 0.00191176
R2429 iovss.n92 iovss.n76 0.00191176
R2430 iovss.n92 iovss.n91 0.00191176
R2431 iovss.n91 iovss.n84 0.00191176
R2432 sg13g2_RCClampResistor_0.pin2.n0 sg13g2_RCClampResistor_0.pin2.t1 10.5567
R2433 sg13g2_RCClampResistor_0.pin2.n0 sg13g2_RCClampResistor_0.pin2.t2 10.286
R2434 sg13g2_RCClampResistor_0.pin2.n1 sg13g2_RCClampResistor_0.pin2.t0 5.0005
R2435 sg13g2_RCClampResistor_0.pin2.n1 sg13g2_RCClampResistor_0.pin2 3.73153
R2436 sg13g2_RCClampResistor_0.pin2 sg13g2_RCClampResistor_0.pin2.n1 0.0214524
R2437 sg13g2_RCClampResistor_0.pin2 sg13g2_RCClampResistor_0.pin2.n0 0.00107971
R2438 vdd.n74 vdd.n73 1.50539
R2439 vdd.n1 vdd.n0 1.5005
R2440 vdd.n69 vdd.n68 1.5005
R2441 vdd.n67 vdd.n66 1.5005
R2442 vdd.n5 vdd.n4 1.5005
R2443 vdd.n61 vdd.n60 1.5005
R2444 vdd.n59 vdd.n58 1.5005
R2445 vdd.n9 vdd.n8 1.5005
R2446 vdd.n53 vdd.n52 1.5005
R2447 vdd.n51 vdd.n50 1.5005
R2448 vdd.n13 vdd.n12 1.5005
R2449 vdd.n45 vdd.n44 1.5005
R2450 vdd.n43 vdd.n42 1.5005
R2451 vdd.n17 vdd.n16 1.5005
R2452 vdd.n37 vdd.n36 1.5005
R2453 vdd.n35 vdd.n34 1.5005
R2454 vdd.n21 vdd.n20 1.5005
R2455 vdd.n29 vdd.n28 1.5005
R2456 vdd.n27 vdd.n26 1.5005
R2457 vdd.n75 vdd 0.6957
R2458 vdd.n73 vdd.n72 0.314786
R2459 vdd.n71 vdd.n70 0.314786
R2460 vdd.n3 vdd.n2 0.314786
R2461 vdd.n65 vdd.n64 0.314786
R2462 vdd.n63 vdd.n62 0.314786
R2463 vdd.n7 vdd.n6 0.314786
R2464 vdd.n57 vdd.n56 0.314786
R2465 vdd.n55 vdd.n54 0.314786
R2466 vdd.n11 vdd.n10 0.314786
R2467 vdd.n49 vdd.n48 0.314786
R2468 vdd.n47 vdd.n46 0.314786
R2469 vdd.n15 vdd.n14 0.314786
R2470 vdd.n41 vdd.n40 0.314786
R2471 vdd.n39 vdd.n38 0.314786
R2472 vdd.n19 vdd.n18 0.314786
R2473 vdd.n33 vdd.n32 0.314786
R2474 vdd.n31 vdd.n30 0.314786
R2475 vdd.n23 vdd.n22 0.314786
R2476 vdd.n24 vdd 0.217715
R2477 vdd.n51 vdd 0.195018
R2478 vdd.n25 vdd.n24 0.146103
R2479 vdd.n26 vdd.n25 0.0354467
R2480 vdd.n25 vdd.n22 0.0314255
R2481 vdd.n28 vdd.n27 0.00921287
R2482 vdd.n28 vdd.n20 0.00921287
R2483 vdd.n35 vdd.n20 0.00921287
R2484 vdd.n36 vdd.n35 0.00921287
R2485 vdd.n36 vdd.n16 0.00921287
R2486 vdd.n43 vdd.n16 0.00921287
R2487 vdd.n44 vdd.n43 0.00921287
R2488 vdd.n44 vdd.n12 0.00921287
R2489 vdd.n51 vdd.n12 0.00921287
R2490 vdd.n52 vdd.n51 0.00921287
R2491 vdd.n52 vdd.n8 0.00921287
R2492 vdd.n59 vdd.n8 0.00921287
R2493 vdd.n60 vdd.n59 0.00921287
R2494 vdd.n60 vdd.n4 0.00921287
R2495 vdd.n67 vdd.n4 0.00921287
R2496 vdd.n68 vdd.n67 0.00921287
R2497 vdd.n68 vdd.n0 0.00921287
R2498 vdd.n74 vdd.n0 0.00921287
R2499 vdd.n26 vdd.n23 0.00538889
R2500 vdd.n29 vdd.n23 0.00538889
R2501 vdd.n30 vdd.n29 0.00538889
R2502 vdd.n30 vdd.n21 0.00538889
R2503 vdd.n33 vdd.n21 0.00538889
R2504 vdd.n34 vdd.n33 0.00538889
R2505 vdd.n34 vdd.n19 0.00538889
R2506 vdd.n37 vdd.n19 0.00538889
R2507 vdd.n38 vdd.n37 0.00538889
R2508 vdd.n38 vdd.n17 0.00538889
R2509 vdd.n41 vdd.n17 0.00538889
R2510 vdd.n42 vdd.n41 0.00538889
R2511 vdd.n42 vdd.n15 0.00538889
R2512 vdd.n45 vdd.n15 0.00538889
R2513 vdd.n46 vdd.n45 0.00538889
R2514 vdd.n46 vdd.n13 0.00538889
R2515 vdd.n49 vdd.n13 0.00538889
R2516 vdd.n50 vdd.n49 0.00538889
R2517 vdd.n50 vdd.n11 0.00538889
R2518 vdd.n53 vdd.n11 0.00538889
R2519 vdd.n54 vdd.n53 0.00538889
R2520 vdd.n54 vdd.n9 0.00538889
R2521 vdd.n57 vdd.n9 0.00538889
R2522 vdd.n58 vdd.n57 0.00538889
R2523 vdd.n58 vdd.n7 0.00538889
R2524 vdd.n61 vdd.n7 0.00538889
R2525 vdd.n62 vdd.n61 0.00538889
R2526 vdd.n62 vdd.n5 0.00538889
R2527 vdd.n65 vdd.n5 0.00538889
R2528 vdd.n66 vdd.n65 0.00538889
R2529 vdd.n66 vdd.n3 0.00538889
R2530 vdd.n69 vdd.n3 0.00538889
R2531 vdd.n70 vdd.n69 0.00538889
R2532 vdd.n70 vdd.n1 0.00538889
R2533 vdd.n73 vdd.n1 0.00538889
R2534 vdd.n27 vdd.n24 0.00485644
R2535 vdd.n75 vdd.n74 0.00485644
R2536 vdd vdd.n75 0.00485644
R2537 vdd.n72 vdd 0.0035
R2538 vdd.n31 vdd.n22 0.0025
R2539 vdd.n32 vdd.n31 0.0025
R2540 vdd.n32 vdd.n18 0.0025
R2541 vdd.n39 vdd.n18 0.0025
R2542 vdd.n40 vdd.n39 0.0025
R2543 vdd.n40 vdd.n14 0.0025
R2544 vdd.n47 vdd.n14 0.0025
R2545 vdd.n48 vdd.n47 0.0025
R2546 vdd.n48 vdd.n10 0.0025
R2547 vdd.n55 vdd.n10 0.0025
R2548 vdd.n56 vdd.n55 0.0025
R2549 vdd.n56 vdd.n6 0.0025
R2550 vdd.n63 vdd.n6 0.0025
R2551 vdd.n64 vdd.n63 0.0025
R2552 vdd.n64 vdd.n2 0.0025
R2553 vdd.n71 vdd.n2 0.0025
R2554 vdd.n72 vdd.n71 0.0025
C0 a_11365_7542# a_11035_7542# 0.37213f
C1 a_4105_7542# a_4435_7542# 0.37213f
C2 a_8065_7542# a_8395_7542# 0.37213f
C3 a_6415_7542# a_6745_7542# 0.37213f
C4 a_5425_7542# a_5755_7542# 0.37213f
C5 a_8725_7542# a_9055_7542# 0.37213f
C6 a_10705_7542# a_10375_7542# 0.37213f
C7 a_5095_7542# a_4765_7542# 0.37213f
C8 iovdd sg13g2_RCClampResistor_0.pin2 90.4337f
C9 a_6085_7542# a_5755_7542# 0.37213f
C10 a_4435_7542# a_4765_7542# 0.37213f
C11 a_3775_7542# a_4105_7542# 0.37213f
C12 a_11695_7542# a_12025_7542# 0.37213f
C13 a_8725_7542# a_8395_7542# 0.37213f
C14 a_7075_7542# a_7405_7542# 0.37213f
C15 a_7405_7542# a_7735_7542# 0.37213f
C16 sg13g2_Clamp_N43N43D4R_0.gate sg13g2_RCClampResistor_0.pin2 21.6731f
C17 a_7075_7542# a_6745_7542# 0.37213f
C18 a_6085_7542# a_6415_7542# 0.37213f
C19 a_10705_7542# a_11035_7542# 0.37213f
C20 a_10045_7542# a_10375_7542# 0.37213f
C21 a_9715_7542# a_10045_7542# 0.37213f
C22 a_9385_7542# a_9055_7542# 0.37213f
C23 a_9385_7542# a_9715_7542# 0.37213f
C24 a_11365_7542# a_11695_7542# 0.37213f
C25 iovdd sg13g2_Clamp_N43N43D4R_0.gate 0.13605p
C26 a_8065_7542# a_7735_7542# 0.37213f
C27 a_5425_7542# a_5095_7542# 0.37213f
C28 iovdd iovss 0.28124p
C29 vdd iovss 0.24621p
C30 a_12025_7542# iovss 3.53966f $ **FLOATING
C31 a_11695_7456# iovss 0.45487f
C32 a_11695_7542# iovss 3.04229f $ **FLOATING
C33 a_11365_7542# iovss 3.04218f $ **FLOATING
C34 a_11365_11542# iovss 0.41716f
C35 a_11035_7456# iovss 0.43382f
C36 a_11035_7542# iovss 3.04229f $ **FLOATING
C37 a_10705_7542# iovss 3.04218f $ **FLOATING
C38 a_10705_11542# iovss 0.41716f
C39 a_10375_7456# iovss 0.43383f
C40 a_10375_7542# iovss 3.04226f $ **FLOATING
C41 a_10045_7542# iovss 3.04218f $ **FLOATING
C42 a_10045_11542# iovss 0.41716f
C43 a_9715_7456# iovss 0.43386f
C44 a_9715_7542# iovss 3.04218f $ **FLOATING
C45 a_9385_7542# iovss 3.04218f $ **FLOATING
C46 a_9385_11542# iovss 0.41716f
C47 a_9055_7456# iovss 0.43385f
C48 a_9055_7542# iovss 3.04218f $ **FLOATING
C49 a_8725_7542# iovss 3.04229f $ **FLOATING
C50 a_8725_11542# iovss 0.41716f
C51 a_8395_7456# iovss 0.43382f
C52 a_8395_7542# iovss 3.04218f $ **FLOATING
C53 a_8065_7542# iovss 3.04229f $ **FLOATING
C54 a_8065_11542# iovss 0.41716f
C55 a_7735_7456# iovss 0.43382f
C56 a_7735_7542# iovss 3.04218f $ **FLOATING
C57 a_7405_7542# iovss 3.04229f $ **FLOATING
C58 a_7405_11542# iovss 0.41716f
C59 a_7075_7456# iovss 0.43384f
C60 a_7075_7542# iovss 3.04218f $ **FLOATING
C61 a_6745_7542# iovss 3.04224f $ **FLOATING
C62 a_6745_11542# iovss 0.41716f
C63 a_6415_7456# iovss 0.43388f
C64 a_6415_7542# iovss 3.04218f $ **FLOATING
C65 a_6085_7542# iovss 3.04218f $ **FLOATING
C66 a_6085_11542# iovss 0.41716f
C67 a_5755_7456# iovss 0.43386f
C68 a_5755_7542# iovss 3.04218f $ **FLOATING
C69 a_5425_7542# iovss 3.04218f $ **FLOATING
C70 a_5425_11542# iovss 0.41716f
C71 a_5095_7456# iovss 0.43386f
C72 a_5095_7542# iovss 3.04229f $ **FLOATING
C73 a_4765_7542# iovss 3.04218f $ **FLOATING
C74 a_4765_11542# iovss 0.41716f
C75 a_4435_7456# iovss 0.43382f
C76 a_4435_7542# iovss 3.04229f $ **FLOATING
C77 a_4105_7542# iovss 3.04218f $ **FLOATING
C78 a_4105_11542# iovss 0.41716f
C79 a_3775_7456# iovss 0.45486f
C80 a_3775_7542# iovss 3.53976f $ **FLOATING
C81 sg13g2_Clamp_N43N43D4R_0.gate iovss 0.2448p
C82 sg13g2_RCClampResistor_0.pin2 iovss 0.20743p
C83 sg13g2_RCClampResistor_0.pin2.t2 iovss 70.6711f
C84 sg13g2_RCClampResistor_0.pin2.t1 iovss 11.3396f
C85 sg13g2_RCClampResistor_0.pin2.n0 iovss 26.362f
C86 sg13g2_RCClampResistor_0.pin2.n1 iovss 0.27407f
C87 iovdd.n0 iovss 0.36472f
C88 iovdd.n1 iovss 0.41335f
C89 iovdd.n2 iovss 0.20667f
C90 iovdd.n3 iovss 0.41335f
C91 iovdd.n4 iovss 0.41335f
C92 iovdd.n5 iovss 0.41335f
C93 iovdd.n6 iovss 0.20667f
C94 iovdd.n7 iovss 0.41335f
C95 iovdd.n8 iovss 0.36472f
C96 iovdd.n9 iovss 0.41335f
C97 iovdd.n10 iovss 0.20667f
C98 iovdd.n11 iovss 0.20667f
C99 iovdd.n12 iovss 0.41335f
C100 iovdd.n13 iovss 0.41335f
C101 iovdd.n14 iovss 0.41335f
C102 iovdd.n15 iovss 0.20667f
C103 iovdd.n16 iovss 0.41335f
C104 iovdd.n17 iovss 0.55377f
C105 iovdd.n18 iovss 5.28752f
C106 iovdd.n19 iovss 0.36472f
C107 iovdd.n20 iovss 0.41335f
C108 iovdd.n21 iovss 0.20667f
C109 iovdd.n22 iovss 0.20667f
C110 iovdd.n23 iovss 0.41335f
C111 iovdd.n24 iovss 0.41335f
C112 iovdd.n25 iovss 0.41335f
C113 iovdd.n26 iovss 0.20667f
C114 iovdd.n27 iovss 0.41335f
C115 iovdd.n28 iovss 0.36472f
C116 iovdd.n29 iovss 0.41335f
C117 iovdd.n30 iovss 0.20667f
C118 iovdd.n31 iovss 0.20667f
C119 iovdd.n32 iovss 0.41335f
C120 iovdd.n33 iovss 0.41335f
C121 iovdd.n34 iovss 0.41335f
C122 iovdd.n35 iovss 0.20667f
C123 iovdd.n36 iovss 0.41335f
C124 iovdd.n37 iovss 0.36472f
C125 iovdd.n38 iovss 0.41335f
C126 iovdd.n39 iovss 0.20667f
C127 iovdd.n40 iovss 0.20667f
C128 iovdd.n41 iovss 0.41335f
C129 iovdd.n42 iovss 0.41335f
C130 iovdd.n43 iovss 0.41335f
C131 iovdd.n44 iovss 0.20667f
C132 iovdd.n45 iovss 0.41335f
C133 iovdd.n46 iovss 5.57115f
C134 iovdd.n47 iovss 0.55377f
C135 iovdd.n48 iovss 0.36472f
C136 iovdd.n49 iovss 0.41335f
C137 iovdd.n50 iovss 0.20667f
C138 iovdd.n51 iovss 0.20667f
C139 iovdd.n52 iovss 0.41335f
C140 iovdd.n53 iovss 0.41335f
C141 iovdd.n54 iovss 0.41335f
C142 iovdd.n55 iovss 0.20667f
C143 iovdd.n56 iovss 0.41335f
C144 iovdd.n57 iovss 0.36472f
C145 iovdd.n58 iovss 0.41335f
C146 iovdd.n59 iovss 0.20667f
C147 iovdd.n60 iovss 0.20667f
C148 iovdd.n61 iovss 0.41335f
C149 iovdd.n62 iovss 0.41335f
C150 iovdd.n63 iovss 0.41335f
C151 iovdd.n64 iovss 0.20667f
C152 iovdd.n65 iovss 0.41335f
C153 iovdd.n66 iovss 0.36472f
C154 iovdd.n67 iovss 0.41335f
C155 iovdd.n68 iovss 0.20667f
C156 iovdd.n69 iovss 0.20667f
C157 iovdd.n70 iovss 0.41335f
C158 iovdd.n71 iovss 0.41335f
C159 iovdd.n72 iovss 0.41335f
C160 iovdd.n73 iovss 0.20667f
C161 iovdd.n74 iovss 0.41335f
C162 iovdd.n75 iovss 0.72898f
C163 iovdd.n76 iovss 1.09416f
C164 iovdd.n137 iovss 0.3215f
C165 iovdd.n138 iovss 0.37437f
C166 iovdd.n149 iovss 1.01796f
C167 iovdd.n150 iovss 1.09416f
C168 iovdd.n590 iovss 1.09416f
C169 iovdd.n591 iovss 1.09416f
C170 iovdd.n592 iovss 0.68385f
C171 iovdd.n606 iovss 5.91164f
C172 iovdd.n625 iovss 0.11636f
C173 iovdd.n667 iovss 13.9526f
C174 iovdd.n668 iovss 1.04766f
C175 iovdd.n669 iovss 1.09416f
C176 iovdd.n673 iovss 0.91225f
C177 iovdd.n674 iovss 0.33417f
C178 iovdd.n675 iovss 0.36472f
C179 iovdd.n676 iovss 0.41335f
C180 iovdd.n677 iovss 0.41335f
C181 iovdd.n678 iovss 0.20667f
C182 iovdd.n679 iovss 0.20667f
C183 iovdd.n680 iovss 0.41335f
C184 iovdd.n681 iovss 0.41335f
C185 iovdd.n682 iovss 0.41335f
C186 iovdd.n683 iovss 0.20667f
C187 iovdd.n684 iovss 0.41335f
C188 iovdd.n685 iovss 1.43358f
C189 iovdd.n686 iovss 0.41335f
C190 iovdd.n687 iovss 0.20667f
C191 iovdd.n688 iovss 0.20667f
C192 iovdd.n689 iovss 0.41335f
C193 iovdd.n690 iovss 0.67757f
C194 iovdd.n691 iovss 0.41335f
C195 iovdd.n692 iovss 0.20667f
C196 iovdd.n693 iovss 0.72924f
C197 iovdd.n694 iovss 0.847f
C198 iovdd.n695 iovss 0.41335f
C199 iovdd.n696 iovss 0.20667f
C200 iovdd.n697 iovss 0.20667f
C201 iovdd.n698 iovss 0.20667f
C202 iovdd.n699 iovss 0.41335f
C203 iovdd.n700 iovss 2.84866f
C204 iovdd.n701 iovss 0.41335f
C205 iovdd.n702 iovss 0.41335f
C206 iovdd.n703 iovss 0.41335f
C207 iovdd.n704 iovss 0.20667f
C208 iovdd.n705 iovss 0.20667f
C209 iovdd.n706 iovss 0.41335f
C210 iovdd.n707 iovss 0.36472f
C211 iovdd.n708 iovss 0.36472f
C212 iovdd.n709 iovss 0.36472f
C213 iovdd.n710 iovss 0.41335f
C214 iovdd.n711 iovss 0.20667f
C215 iovdd.n712 iovss 0.20667f
C216 iovdd.n713 iovss 0.20667f
C217 iovdd.n714 iovss 0.41335f
C218 iovdd.n715 iovss 0.41335f
C219 iovdd.n716 iovss 0.41335f
C220 iovdd.n717 iovss 0.41335f
C221 iovdd.n718 iovss 0.41335f
C222 iovdd.n719 iovss 0.41335f
C223 iovdd.n720 iovss 0.20667f
C224 iovdd.n721 iovss 0.41335f
C225 iovdd.n722 iovss 0.36472f
C226 iovdd.n723 iovss 0.41335f
C227 iovdd.n724 iovss 0.20667f
C228 iovdd.n725 iovss 0.20667f
C229 iovdd.n726 iovss 0.20667f
C230 iovdd.n727 iovss 0.41335f
C231 iovdd.n728 iovss 0.41335f
C232 iovdd.n729 iovss 0.41335f
C233 iovdd.n730 iovss 0.41335f
C234 iovdd.n731 iovss 0.41335f
C235 iovdd.n732 iovss 0.41335f
C236 iovdd.n733 iovss 0.20667f
C237 iovdd.n734 iovss 0.41335f
C238 iovdd.n735 iovss 0.36472f
C239 iovdd.n736 iovss 0.41335f
C240 iovdd.n737 iovss 0.20667f
C241 iovdd.n738 iovss 0.20667f
C242 iovdd.n739 iovss 0.20667f
C243 iovdd.n740 iovss 0.41335f
C244 iovdd.n741 iovss 0.41335f
C245 iovdd.n742 iovss 0.41335f
C246 iovdd.n743 iovss 0.41335f
C247 iovdd.n744 iovss 0.41335f
C248 iovdd.n745 iovss 0.41335f
C249 iovdd.n746 iovss 0.20667f
C250 iovdd.n747 iovss 0.41335f
C251 iovdd.n748 iovss 0.20667f
C252 iovdd.n749 iovss 0.41335f
C253 iovdd.t89 iovss 4.85281f
C254 iovdd.n804 iovss 0.31833f
C255 iovdd.n807 iovss 0.46925f
C256 iovdd.n808 iovss 0.41335f
C257 iovdd.n809 iovss 0.41335f
C258 iovdd.n810 iovss 0.20667f
C259 iovdd.n811 iovss 0.41335f
C260 iovdd.n812 iovss 0.27308f
C261 iovdd.n813 iovss 0.36472f
C262 iovdd.n814 iovss 0.41335f
C263 iovdd.n815 iovss 0.20667f
C264 iovdd.n816 iovss 0.20667f
C265 iovdd.n817 iovss 0.20667f
C266 iovdd.n818 iovss 0.41335f
C267 iovdd.n819 iovss 0.41335f
C268 iovdd.n820 iovss 0.41335f
C269 iovdd.n821 iovss 0.41335f
C270 iovdd.n822 iovss 0.41335f
C271 iovdd.n823 iovss 0.41335f
C272 iovdd.n824 iovss 0.20667f
C273 iovdd.n825 iovss 0.41335f
C274 iovdd.n826 iovss 0.36472f
C275 iovdd.n827 iovss 0.41335f
C276 iovdd.n828 iovss 0.20667f
C277 iovdd.n829 iovss 0.20667f
C278 iovdd.n830 iovss 0.20667f
C279 iovdd.n831 iovss 0.41335f
C280 iovdd.n832 iovss 0.41335f
C281 iovdd.n833 iovss 0.41335f
C282 iovdd.n834 iovss 0.41335f
C283 iovdd.n835 iovss 0.41335f
C284 iovdd.n836 iovss 0.41335f
C285 iovdd.n837 iovss 0.20667f
C286 iovdd.n838 iovss 0.41335f
C287 iovdd.n839 iovss 0.41335f
C288 iovdd.n840 iovss 0.20667f
C289 iovdd.n841 iovss 0.20667f
C290 iovdd.n842 iovss 0.20667f
C291 iovdd.n843 iovss 0.41335f
C292 iovdd.n844 iovss 0.41335f
C293 iovdd.n845 iovss 0.41335f
C294 iovdd.n846 iovss 0.41335f
C295 iovdd.n847 iovss 0.41335f
C296 iovdd.n848 iovss 0.41335f
C297 iovdd.n849 iovss 0.20667f
C298 iovdd.n850 iovss 0.41335f
C299 iovdd.n851 iovss 0.33417f
C300 iovdd.n852 iovss 0.36472f
C301 iovdd.n853 iovss 0.41335f
C302 iovdd.n854 iovss 0.20667f
C303 iovdd.n855 iovss 0.20667f
C304 iovdd.n856 iovss 0.20667f
C305 iovdd.n857 iovss 0.41335f
C306 iovdd.n858 iovss 0.41335f
C307 iovdd.n859 iovss 0.41335f
C308 iovdd.n860 iovss 0.41335f
C309 iovdd.n861 iovss 0.41335f
C310 iovdd.n862 iovss 0.41335f
C311 iovdd.n863 iovss 0.20667f
C312 iovdd.n864 iovss 0.41335f
C313 iovdd.n865 iovss 0.41335f
C314 iovdd.n866 iovss 0.62219f
C315 iovdd.n867 iovss 0.72119f
C316 iovdd.n868 iovss 0.8267f
C317 iovdd.n869 iovss 0.4559f
C318 iovdd.n870 iovss 0.36472f
C319 iovdd.n871 iovss 0.41335f
C320 iovdd.n872 iovss 0.20667f
C321 iovdd.n873 iovss 0.20667f
C322 iovdd.n874 iovss 0.41335f
C323 iovdd.n875 iovss 0.41335f
C324 iovdd.n876 iovss 0.20667f
C325 iovdd.n877 iovss 0.20667f
C326 iovdd.n878 iovss 0.41335f
C327 iovdd.n879 iovss 0.36472f
C328 iovdd.n880 iovss 0.36472f
C329 iovdd.n881 iovss 0.36472f
C330 iovdd.n882 iovss 0.41335f
C331 iovdd.n883 iovss 0.20667f
C332 iovdd.n884 iovss 0.20667f
C333 iovdd.n885 iovss 0.41335f
C334 iovdd.n886 iovss 0.41335f
C335 iovdd.n887 iovss 0.20667f
C336 iovdd.n888 iovss 0.20667f
C337 iovdd.n889 iovss 0.41335f
C338 iovdd.n890 iovss 0.21291f
C339 iovdd.n891 iovss 0.36472f
C340 iovdd.n892 iovss 0.36472f
C341 iovdd.n893 iovss 0.41335f
C342 iovdd.n894 iovss 0.20667f
C343 iovdd.n895 iovss 0.20667f
C344 iovdd.n896 iovss 0.41335f
C345 iovdd.n897 iovss 0.41335f
C346 iovdd.n898 iovss 0.20667f
C347 iovdd.n899 iovss 0.20667f
C348 iovdd.n900 iovss 0.41335f
C349 iovdd.n901 iovss 0.36472f
C350 iovdd.n902 iovss 0.36472f
C351 iovdd.n903 iovss 0.36472f
C352 iovdd.n904 iovss 0.41335f
C353 iovdd.n905 iovss 0.20667f
C354 iovdd.n906 iovss 0.20667f
C355 iovdd.n907 iovss 0.41335f
C356 iovdd.n908 iovss 0.41335f
C357 iovdd.n909 iovss 0.20667f
C358 iovdd.n910 iovss 0.20667f
C359 iovdd.n911 iovss 0.41335f
C360 iovdd.n912 iovss 0.36472f
C361 iovdd.n913 iovss 0.36472f
C362 iovdd.n914 iovss 0.36472f
C363 iovdd.n915 iovss 0.41335f
C364 iovdd.n916 iovss 0.20667f
C365 iovdd.n917 iovss 0.20667f
C366 iovdd.n918 iovss 0.41335f
C367 iovdd.n919 iovss 0.41335f
C368 iovdd.n920 iovss 0.20667f
C369 iovdd.n921 iovss 0.20667f
C370 iovdd.n922 iovss 0.41335f
C371 iovdd.n923 iovss 0.27399f
C372 iovdd.n924 iovss 0.36472f
C373 iovdd.n925 iovss 0.41335f
C374 iovdd.n926 iovss 0.20667f
C375 iovdd.n927 iovss 0.20667f
C376 iovdd.n928 iovss 0.41335f
C377 iovdd.n929 iovss 0.41335f
C378 iovdd.n930 iovss 0.20667f
C379 iovdd.n931 iovss 0.20667f
C380 iovdd.n932 iovss 0.41335f
C381 iovdd.n933 iovss 0.36472f
C382 iovdd.n934 iovss 0.36472f
C383 iovdd.n935 iovss 0.36472f
C384 iovdd.n936 iovss 0.41335f
C385 iovdd.n937 iovss 0.20667f
C386 iovdd.n938 iovss 0.20667f
C387 iovdd.n939 iovss 0.41335f
C388 iovdd.n940 iovss 0.41335f
C389 iovdd.n941 iovss 0.20667f
C390 iovdd.n942 iovss 0.20667f
C391 iovdd.n943 iovss 0.41335f
C392 iovdd.n944 iovss 0.36472f
C393 iovdd.n945 iovss 0.36472f
C394 iovdd.n946 iovss 0.36472f
C395 iovdd.n947 iovss 0.41335f
C396 iovdd.n948 iovss 0.20667f
C397 iovdd.n949 iovss 0.20667f
C398 iovdd.n950 iovss 0.41335f
C399 iovdd.n951 iovss 0.41335f
C400 iovdd.n952 iovss 0.20667f
C401 iovdd.n953 iovss 0.20667f
C402 iovdd.n954 iovss 0.41335f
C403 iovdd.n955 iovss 0.21291f
C404 iovdd.n956 iovss 0.55377f
C405 iovdd.n957 iovss 0.36472f
C406 iovdd.n958 iovss 0.41335f
C407 iovdd.n959 iovss 0.20667f
C408 iovdd.n960 iovss 0.20667f
C409 iovdd.n961 iovss 0.41335f
C410 iovdd.n962 iovss 0.41335f
C411 iovdd.n963 iovss 0.41335f
C412 iovdd.n964 iovss 0.20667f
C413 iovdd.n965 iovss 0.41335f
C414 iovdd.n966 iovss 0.72918f
C415 iovdd.n967 iovss 0.20667f
C416 iovdd.n968 iovss 0.20667f
C417 iovdd.n969 iovss 0.41335f
C418 iovdd.n970 iovss 0.64142f
C419 iovdd.n971 iovss 1.4245f
C420 iovdd.n972 iovss 0.41335f
C421 iovdd.n973 iovss 0.20667f
C422 iovdd.n974 iovss 0.20667f
C423 iovdd.n975 iovss 0.41335f
C424 iovdd.n976 iovss 0.847f
C425 iovdd.n977 iovss 1.43358f
C426 iovdd.n978 iovss 0.36472f
C427 iovdd.n979 iovss 0.41335f
C428 iovdd.n980 iovss 0.20667f
C429 iovdd.n981 iovss 0.20667f
C430 iovdd.n982 iovss 0.20667f
C431 iovdd.n983 iovss 0.41335f
C432 iovdd.n984 iovss 0.41335f
C433 iovdd.n985 iovss 0.41335f
C434 iovdd.n986 iovss 0.41335f
C435 iovdd.n987 iovss 0.41335f
C436 iovdd.n988 iovss 0.20667f
C437 iovdd.n989 iovss 0.20667f
C438 iovdd.n990 iovss 0.41335f
C439 iovdd.n991 iovss 0.36472f
C440 iovdd.n992 iovss 0.33417f
C441 iovdd.n993 iovss 1.10084f
C442 iovdd.n994 iovss 0.21291f
C443 iovdd.n995 iovss 0.41335f
C444 iovdd.n996 iovss 0.20667f
C445 iovdd.n997 iovss 0.20667f
C446 iovdd.n998 iovss 0.20667f
C447 iovdd.n999 iovss 0.41335f
C448 iovdd.n1000 iovss 0.41335f
C449 iovdd.n1001 iovss 0.41335f
C450 iovdd.n1002 iovss 0.41335f
C451 iovdd.n1003 iovss 0.41335f
C452 iovdd.n1004 iovss 0.20667f
C453 iovdd.n1005 iovss 0.20667f
C454 iovdd.n1006 iovss 0.41335f
C455 iovdd.n1007 iovss 0.36472f
C456 iovdd.n1008 iovss 0.36472f
C457 iovdd.n1009 iovss 0.36472f
C458 iovdd.n1010 iovss 0.41335f
C459 iovdd.n1011 iovss 0.20667f
C460 iovdd.n1012 iovss 0.20667f
C461 iovdd.n1013 iovss 0.20667f
C462 iovdd.n1014 iovss 0.41335f
C463 iovdd.n1015 iovss 0.41335f
C464 iovdd.n1016 iovss 0.41335f
C465 iovdd.n1017 iovss 0.41335f
C466 iovdd.n1018 iovss 0.41335f
C467 iovdd.n1019 iovss 0.20667f
C468 iovdd.n1020 iovss 0.20667f
C469 iovdd.n1021 iovss 0.41335f
C470 iovdd.n1022 iovss 0.36472f
C471 iovdd.n1023 iovss 0.36472f
C472 iovdd.n1024 iovss 0.36472f
C473 iovdd.n1025 iovss 0.41335f
C474 iovdd.n1026 iovss 0.20667f
C475 iovdd.n1027 iovss 0.20667f
C476 iovdd.n1028 iovss 0.20667f
C477 iovdd.n1029 iovss 0.41335f
C478 iovdd.n1030 iovss 0.41335f
C479 iovdd.n1031 iovss 0.41335f
C480 iovdd.n1032 iovss 0.41335f
C481 iovdd.n1033 iovss 0.41335f
C482 iovdd.n1034 iovss 0.20667f
C483 iovdd.n1035 iovss 0.20667f
C484 iovdd.n1036 iovss 0.41335f
C485 iovdd.n1037 iovss 0.36472f
C486 iovdd.n1038 iovss 0.27399f
C487 iovdd.n1039 iovss 5.45632f
C488 iovdd.n1040 iovss 0.27308f
C489 iovdd.n1041 iovss 0.41335f
C490 iovdd.n1042 iovss 0.20667f
C491 iovdd.n1043 iovss 0.20667f
C492 iovdd.n1044 iovss 0.20667f
C493 iovdd.n1045 iovss 0.41335f
C494 iovdd.n1046 iovss 0.41335f
C495 iovdd.n1047 iovss 0.41335f
C496 iovdd.n1048 iovss 0.41335f
C497 iovdd.n1049 iovss 0.41335f
C498 iovdd.n1050 iovss 0.20667f
C499 iovdd.n1051 iovss 0.20667f
C500 iovdd.n1052 iovss 0.41335f
C501 iovdd.n1053 iovss 0.36472f
C502 iovdd.n1054 iovss 0.36472f
C503 iovdd.n1055 iovss 0.36472f
C504 iovdd.n1056 iovss 0.41335f
C505 iovdd.n1057 iovss 0.20667f
C506 iovdd.n1058 iovss 0.20667f
C507 iovdd.n1059 iovss 0.20667f
C508 iovdd.n1060 iovss 0.41335f
C509 iovdd.n1061 iovss 0.41335f
C510 iovdd.n1062 iovss 0.41335f
C511 iovdd.n1063 iovss 0.41335f
C512 iovdd.n1064 iovss 0.41335f
C513 iovdd.n1065 iovss 0.20667f
C514 iovdd.n1066 iovss 0.20667f
C515 iovdd.n1067 iovss 0.41335f
C516 iovdd.n1068 iovss 0.36472f
C517 iovdd.n1069 iovss 0.36472f
C518 iovdd.n1070 iovss 0.36472f
C519 iovdd.n1071 iovss 0.41335f
C520 iovdd.n1072 iovss 0.20667f
C521 iovdd.n1073 iovss 0.20667f
C522 iovdd.n1074 iovss 0.20667f
C523 iovdd.n1075 iovss 0.41335f
C524 iovdd.n1076 iovss 0.41335f
C525 iovdd.n1077 iovss 0.41335f
C526 iovdd.n1078 iovss 0.41335f
C527 iovdd.n1079 iovss 0.41335f
C528 iovdd.n1080 iovss 0.20667f
C529 iovdd.n1081 iovss 0.20667f
C530 iovdd.n1082 iovss 0.41335f
C531 iovdd.n1083 iovss 0.36472f
C532 iovdd.n1084 iovss 0.21291f
C533 iovdd.n1085 iovss 5.45632f
C534 iovdd.n1086 iovss 0.33417f
C535 iovdd.n1087 iovss 0.41335f
C536 iovdd.n1088 iovss 0.20667f
C537 iovdd.n1089 iovss 0.20667f
C538 iovdd.n1090 iovss 0.20667f
C539 iovdd.n1091 iovss 0.41335f
C540 iovdd.n1092 iovss 0.41335f
C541 iovdd.n1093 iovss 0.41335f
C542 iovdd.n1094 iovss 0.41335f
C543 iovdd.n1095 iovss 0.41335f
C544 iovdd.n1096 iovss 0.20667f
C545 iovdd.n1097 iovss 0.20667f
C546 iovdd.n1098 iovss 0.41335f
C547 iovdd.n1099 iovss 0.36472f
C548 iovdd.n1100 iovss 0.36472f
C549 iovdd.n1101 iovss 0.36472f
C550 iovdd.n1102 iovss 0.41335f
C551 iovdd.n1103 iovss 0.20667f
C552 iovdd.n1104 iovss 0.20667f
C553 iovdd.n1105 iovss 0.20667f
C554 iovdd.n1106 iovss 0.41335f
C555 iovdd.n1107 iovss 1.4245f
C556 iovdd.n1108 iovss 0.64142f
C557 iovdd.n1109 iovss 0.72419f
C558 iovdd.n1110 iovss 0.51669f
C559 iovdd.n1111 iovss 0.4559f
C560 sg13g2_Clamp_N43N43D4R_0.gate.t66 iovss 0.9055f
C561 sg13g2_Clamp_N43N43D4R_0.gate.t109 iovss 0.51153f
C562 sg13g2_Clamp_N43N43D4R_0.gate.n0 iovss 0.11866f
C563 sg13g2_Clamp_N43N43D4R_0.gate.t70 iovss 0.9055f
C564 sg13g2_Clamp_N43N43D4R_0.gate.t85 iovss 0.51153f
C565 sg13g2_Clamp_N43N43D4R_0.gate.n2 iovss 0.36603f
C566 sg13g2_Clamp_N43N43D4R_0.gate.t88 iovss 0.9055f
C567 sg13g2_Clamp_N43N43D4R_0.gate.t32 iovss 0.51153f
C568 sg13g2_Clamp_N43N43D4R_0.gate.n4 iovss 0.2025f
C569 sg13g2_Clamp_N43N43D4R_0.gate.t37 iovss 0.9055f
C570 sg13g2_Clamp_N43N43D4R_0.gate.t99 iovss 0.51153f
C571 sg13g2_Clamp_N43N43D4R_0.gate.n6 iovss 0.2025f
C572 sg13g2_Clamp_N43N43D4R_0.gate.t51 iovss 0.9055f
C573 sg13g2_Clamp_N43N43D4R_0.gate.t68 iovss 0.51153f
C574 sg13g2_Clamp_N43N43D4R_0.gate.n8 iovss 0.2025f
C575 sg13g2_Clamp_N43N43D4R_0.gate.t60 iovss 0.9055f
C576 sg13g2_Clamp_N43N43D4R_0.gate.t103 iovss 0.51153f
C577 sg13g2_Clamp_N43N43D4R_0.gate.n10 iovss 0.2025f
C578 sg13g2_Clamp_N43N43D4R_0.gate.t75 iovss 0.9055f
C579 sg13g2_Clamp_N43N43D4R_0.gate.t89 iovss 0.51153f
C580 sg13g2_Clamp_N43N43D4R_0.gate.n12 iovss 0.2025f
C581 sg13g2_Clamp_N43N43D4R_0.gate.t98 iovss 0.9055f
C582 sg13g2_Clamp_N43N43D4R_0.gate.t47 iovss 0.51153f
C583 sg13g2_Clamp_N43N43D4R_0.gate.n14 iovss 0.2025f
C584 sg13g2_Clamp_N43N43D4R_0.gate.t58 iovss 0.9055f
C585 sg13g2_Clamp_N43N43D4R_0.gate.t72 iovss 0.51153f
C586 sg13g2_Clamp_N43N43D4R_0.gate.n16 iovss 0.2025f
C587 sg13g2_Clamp_N43N43D4R_0.gate.t53 iovss 0.9055f
C588 sg13g2_Clamp_N43N43D4R_0.gate.t69 iovss 0.51153f
C589 sg13g2_Clamp_N43N43D4R_0.gate.n18 iovss 0.2025f
C590 sg13g2_Clamp_N43N43D4R_0.gate.t45 iovss 0.9055f
C591 sg13g2_Clamp_N43N43D4R_0.gate.t106 iovss 0.51153f
C592 sg13g2_Clamp_N43N43D4R_0.gate.n20 iovss 0.2025f
C593 sg13g2_Clamp_N43N43D4R_0.gate.t36 iovss 0.9055f
C594 sg13g2_Clamp_N43N43D4R_0.gate.t50 iovss 0.51153f
C595 sg13g2_Clamp_N43N43D4R_0.gate.n22 iovss 0.2025f
C596 sg13g2_Clamp_N43N43D4R_0.gate.t67 iovss 0.9055f
C597 sg13g2_Clamp_N43N43D4R_0.gate.t110 iovss 0.51153f
C598 sg13g2_Clamp_N43N43D4R_0.gate.n24 iovss 0.2025f
C599 sg13g2_Clamp_N43N43D4R_0.gate.t56 iovss 0.9055f
C600 sg13g2_Clamp_N43N43D4R_0.gate.t102 iovss 0.51153f
C601 sg13g2_Clamp_N43N43D4R_0.gate.n26 iovss 0.2025f
C602 sg13g2_Clamp_N43N43D4R_0.gate.t33 iovss 0.9055f
C603 sg13g2_Clamp_N43N43D4R_0.gate.t49 iovss 0.51153f
C604 sg13g2_Clamp_N43N43D4R_0.gate.n28 iovss 0.2025f
C605 sg13g2_Clamp_N43N43D4R_0.gate.t34 iovss 0.9055f
C606 sg13g2_Clamp_N43N43D4R_0.gate.t105 iovss 0.51153f
C607 sg13g2_Clamp_N43N43D4R_0.gate.n30 iovss 0.2025f
C608 sg13g2_Clamp_N43N43D4R_0.gate.t86 iovss 0.9055f
C609 sg13g2_Clamp_N43N43D4R_0.gate.t96 iovss 0.51153f
C610 sg13g2_Clamp_N43N43D4R_0.gate.n32 iovss 0.2025f
C611 sg13g2_Clamp_N43N43D4R_0.gate.t41 iovss 0.9055f
C612 sg13g2_Clamp_N43N43D4R_0.gate.t55 iovss 0.51153f
C613 sg13g2_Clamp_N43N43D4R_0.gate.n34 iovss 0.2025f
C614 sg13g2_Clamp_N43N43D4R_0.gate.t65 iovss 0.9055f
C615 sg13g2_Clamp_N43N43D4R_0.gate.t82 iovss 0.51153f
C616 sg13g2_Clamp_N43N43D4R_0.gate.n36 iovss 0.2025f
C617 sg13g2_Clamp_N43N43D4R_0.gate.t62 iovss 0.9055f
C618 sg13g2_Clamp_N43N43D4R_0.gate.t78 iovss 0.51153f
C619 sg13g2_Clamp_N43N43D4R_0.gate.n38 iovss 0.2025f
C620 sg13g2_Clamp_N43N43D4R_0.gate.t54 iovss 0.9055f
C621 sg13g2_Clamp_N43N43D4R_0.gate.t108 iovss 0.51153f
C622 sg13g2_Clamp_N43N43D4R_0.gate.n40 iovss 0.2025f
C623 sg13g2_Clamp_N43N43D4R_0.gate.t46 iovss 0.9055f
C624 sg13g2_Clamp_N43N43D4R_0.gate.t61 iovss 0.51153f
C625 sg13g2_Clamp_N43N43D4R_0.gate.n42 iovss 0.2025f
C626 sg13g2_Clamp_N43N43D4R_0.gate.t77 iovss 0.9055f
C627 sg13g2_Clamp_N43N43D4R_0.gate.t115 iovss 0.51153f
C628 sg13g2_Clamp_N43N43D4R_0.gate.n44 iovss 0.2025f
C629 sg13g2_Clamp_N43N43D4R_0.gate.t31 iovss 0.9055f
C630 sg13g2_Clamp_N43N43D4R_0.gate.t104 iovss 0.51153f
C631 sg13g2_Clamp_N43N43D4R_0.gate.n46 iovss 0.2025f
C632 sg13g2_Clamp_N43N43D4R_0.gate.t42 iovss 0.9055f
C633 sg13g2_Clamp_N43N43D4R_0.gate.t57 iovss 0.51153f
C634 sg13g2_Clamp_N43N43D4R_0.gate.n48 iovss 0.2025f
C635 sg13g2_Clamp_N43N43D4R_0.gate.t48 iovss 0.9055f
C636 sg13g2_Clamp_N43N43D4R_0.gate.t101 iovss 0.51153f
C637 sg13g2_Clamp_N43N43D4R_0.gate.n50 iovss 0.2025f
C638 sg13g2_Clamp_N43N43D4R_0.gate.t63 iovss 0.9055f
C639 sg13g2_Clamp_N43N43D4R_0.gate.t80 iovss 0.51153f
C640 sg13g2_Clamp_N43N43D4R_0.gate.n52 iovss 0.2025f
C641 sg13g2_Clamp_N43N43D4R_0.gate.t90 iovss 0.9055f
C642 sg13g2_Clamp_N43N43D4R_0.gate.t35 iovss 0.51153f
C643 sg13g2_Clamp_N43N43D4R_0.gate.n54 iovss 0.2025f
C644 sg13g2_Clamp_N43N43D4R_0.gate.t87 iovss 0.9055f
C645 sg13g2_Clamp_N43N43D4R_0.gate.t97 iovss 0.51153f
C646 sg13g2_Clamp_N43N43D4R_0.gate.n56 iovss 0.2025f
C647 sg13g2_Clamp_N43N43D4R_0.gate.t43 iovss 0.9055f
C648 sg13g2_Clamp_N43N43D4R_0.gate.t59 iovss 0.51153f
C649 sg13g2_Clamp_N43N43D4R_0.gate.n58 iovss 0.2025f
C650 sg13g2_Clamp_N43N43D4R_0.gate.t74 iovss 0.9055f
C651 sg13g2_Clamp_N43N43D4R_0.gate.t112 iovss 0.51153f
C652 sg13g2_Clamp_N43N43D4R_0.gate.n60 iovss 0.2025f
C653 sg13g2_Clamp_N43N43D4R_0.gate.t92 iovss 0.9055f
C654 sg13g2_Clamp_N43N43D4R_0.gate.t39 iovss 0.51153f
C655 sg13g2_Clamp_N43N43D4R_0.gate.n62 iovss 0.2025f
C656 sg13g2_Clamp_N43N43D4R_0.gate.t93 iovss 0.9055f
C657 sg13g2_Clamp_N43N43D4R_0.gate.t40 iovss 0.51153f
C658 sg13g2_Clamp_N43N43D4R_0.gate.n64 iovss 0.2025f
C659 sg13g2_Clamp_N43N43D4R_0.gate.t44 iovss 0.9055f
C660 sg13g2_Clamp_N43N43D4R_0.gate.t100 iovss 0.51153f
C661 sg13g2_Clamp_N43N43D4R_0.gate.n66 iovss 0.2025f
C662 sg13g2_Clamp_N43N43D4R_0.gate.t79 iovss 0.9055f
C663 sg13g2_Clamp_N43N43D4R_0.gate.t116 iovss 0.51153f
C664 sg13g2_Clamp_N43N43D4R_0.gate.n68 iovss 0.2025f
C665 sg13g2_Clamp_N43N43D4R_0.gate.t83 iovss 0.9055f
C666 sg13g2_Clamp_N43N43D4R_0.gate.t94 iovss 0.51153f
C667 sg13g2_Clamp_N43N43D4R_0.gate.n70 iovss 0.2025f
C668 sg13g2_Clamp_N43N43D4R_0.gate.t84 iovss 0.9055f
C669 sg13g2_Clamp_N43N43D4R_0.gate.t95 iovss 0.51153f
C670 sg13g2_Clamp_N43N43D4R_0.gate.n72 iovss 0.2025f
C671 sg13g2_Clamp_N43N43D4R_0.gate.t71 iovss 0.9055f
C672 sg13g2_Clamp_N43N43D4R_0.gate.t111 iovss 0.51153f
C673 sg13g2_Clamp_N43N43D4R_0.gate.n74 iovss 0.2025f
C674 sg13g2_Clamp_N43N43D4R_0.gate.t64 iovss 0.9055f
C675 sg13g2_Clamp_N43N43D4R_0.gate.t81 iovss 0.51153f
C676 sg13g2_Clamp_N43N43D4R_0.gate.n76 iovss 0.2025f
C677 sg13g2_Clamp_N43N43D4R_0.gate.t91 iovss 0.9055f
C678 sg13g2_Clamp_N43N43D4R_0.gate.t38 iovss 0.51153f
C679 sg13g2_Clamp_N43N43D4R_0.gate.n78 iovss 0.2025f
C680 sg13g2_Clamp_N43N43D4R_0.gate.t52 iovss 0.9055f
C681 sg13g2_Clamp_N43N43D4R_0.gate.t107 iovss 0.51153f
C682 sg13g2_Clamp_N43N43D4R_0.gate.n80 iovss 0.2025f
C683 sg13g2_Clamp_N43N43D4R_0.gate.t73 iovss 0.9055f
C684 sg13g2_Clamp_N43N43D4R_0.gate.t113 iovss 0.51153f
C685 sg13g2_Clamp_N43N43D4R_0.gate.n82 iovss 0.2025f
C686 sg13g2_Clamp_N43N43D4R_0.gate.t76 iovss 0.9055f
C687 sg13g2_Clamp_N43N43D4R_0.gate.t114 iovss 0.51153f
C688 sg13g2_Clamp_N43N43D4R_0.gate.n84 iovss 0.22436f
C689 sg13g2_Clamp_N43N43D4R_0.gate.t24 iovss 0.3917f
C690 sg13g2_Clamp_N43N43D4R_0.gate.t18 iovss 0.38065f
C691 sg13g2_Clamp_N43N43D4R_0.gate.n86 iovss 2.25104f
C692 sg13g2_Clamp_N43N43D4R_0.gate.t19 iovss 0.38065f
C693 sg13g2_Clamp_N43N43D4R_0.gate.n87 iovss 1.42996f
C694 sg13g2_Clamp_N43N43D4R_0.gate.t23 iovss 0.38065f
C695 sg13g2_Clamp_N43N43D4R_0.gate.n88 iovss 1.42996f
C696 sg13g2_Clamp_N43N43D4R_0.gate.t21 iovss 0.38065f
C697 sg13g2_Clamp_N43N43D4R_0.gate.n89 iovss 1.42996f
C698 sg13g2_Clamp_N43N43D4R_0.gate.t20 iovss 0.38065f
C699 sg13g2_Clamp_N43N43D4R_0.gate.n90 iovss 1.42996f
C700 sg13g2_Clamp_N43N43D4R_0.gate.t7 iovss 0.38065f
C701 sg13g2_Clamp_N43N43D4R_0.gate.n91 iovss 1.42996f
C702 sg13g2_Clamp_N43N43D4R_0.gate.t6 iovss 0.38065f
C703 sg13g2_Clamp_N43N43D4R_0.gate.n92 iovss 1.42996f
C704 sg13g2_Clamp_N43N43D4R_0.gate.t3 iovss 0.38065f
C705 sg13g2_Clamp_N43N43D4R_0.gate.n93 iovss 1.42996f
C706 sg13g2_Clamp_N43N43D4R_0.gate.t2 iovss 0.38065f
C707 sg13g2_Clamp_N43N43D4R_0.gate.n94 iovss 1.42996f
C708 sg13g2_Clamp_N43N43D4R_0.gate.t5 iovss 0.38065f
C709 sg13g2_Clamp_N43N43D4R_0.gate.n95 iovss 1.42996f
C710 sg13g2_Clamp_N43N43D4R_0.gate.t4 iovss 0.38065f
C711 sg13g2_Clamp_N43N43D4R_0.gate.n96 iovss 1.42996f
C712 sg13g2_Clamp_N43N43D4R_0.gate.t11 iovss 0.38065f
C713 sg13g2_Clamp_N43N43D4R_0.gate.n97 iovss 1.42996f
C714 sg13g2_Clamp_N43N43D4R_0.gate.t1 iovss 0.38058f
C715 sg13g2_Clamp_N43N43D4R_0.gate.n98 iovss 1.43003f
C716 sg13g2_Clamp_N43N43D4R_0.gate.t0 iovss 0.38065f
C717 sg13g2_Clamp_N43N43D4R_0.gate.n99 iovss 1.42996f
C718 sg13g2_Clamp_N43N43D4R_0.gate.t13 iovss 0.38065f
C719 sg13g2_Clamp_N43N43D4R_0.gate.n100 iovss 1.42996f
C720 sg13g2_Clamp_N43N43D4R_0.gate.t12 iovss 0.38065f
C721 sg13g2_Clamp_N43N43D4R_0.gate.n101 iovss 1.42996f
C722 sg13g2_Clamp_N43N43D4R_0.gate.t17 iovss 0.38065f
C723 sg13g2_Clamp_N43N43D4R_0.gate.n102 iovss 1.42996f
C724 sg13g2_Clamp_N43N43D4R_0.gate.t16 iovss 0.38065f
C725 sg13g2_Clamp_N43N43D4R_0.gate.n103 iovss 1.42996f
C726 sg13g2_Clamp_N43N43D4R_0.gate.t22 iovss 0.38065f
C727 sg13g2_Clamp_N43N43D4R_0.gate.n104 iovss 1.42996f
C728 sg13g2_Clamp_N43N43D4R_0.gate.t15 iovss 0.38065f
C729 sg13g2_Clamp_N43N43D4R_0.gate.n105 iovss 1.42996f
C730 sg13g2_Clamp_N43N43D4R_0.gate.t14 iovss 0.38065f
C731 sg13g2_Clamp_N43N43D4R_0.gate.n106 iovss 1.42996f
C732 sg13g2_Clamp_N43N43D4R_0.gate.t9 iovss 0.38065f
C733 sg13g2_Clamp_N43N43D4R_0.gate.n107 iovss 1.42996f
C734 sg13g2_Clamp_N43N43D4R_0.gate.t8 iovss 0.38065f
C735 sg13g2_Clamp_N43N43D4R_0.gate.n108 iovss 1.42996f
C736 sg13g2_Clamp_N43N43D4R_0.gate.t10 iovss 0.38066f
C737 sg13g2_Clamp_N43N43D4R_0.gate.n109 iovss 12.0539f
C738 sg13g2_Clamp_N43N43D4R_0.gate.t29 iovss 0.5001f
C739 sg13g2_Clamp_N43N43D4R_0.gate.t27 iovss 0.5001f
C740 sg13g2_Clamp_N43N43D4R_0.gate.t25 iovss 0.5001f
C741 sg13g2_Clamp_N43N43D4R_0.gate.n110 iovss 15.0457f
C742 sg13g2_Clamp_N43N43D4R_0.gate.t30 iovss 0.5001f
C743 sg13g2_Clamp_N43N43D4R_0.gate.t28 iovss 0.5001f
C744 sg13g2_Clamp_N43N43D4R_0.gate.t26 iovss 0.5001f
C745 sg13g2_Clamp_N43N43D4R_0.gate.n111 iovss 5.58433f
.ends

