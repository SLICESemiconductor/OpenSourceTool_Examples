* NGSPICE file created from sg13g2_IOPadInOut30mA_flat.ext - technology: ihp-sg13g2

.subckt sg13g2_IOPadInOut30mA_flat p2c c2p_en c2p pad vdd vss iovdd iovss
X0 vdd.t11 a_12038_31490# p2c.t1 vdd.t0 sg13_lv_pmos ad=1.615p pd=10.18u as=1.615p ps=10.18u w=4.75u l=0.13u
X1 sg13g2_GateDecode_0.pgate.t2 iovdd.t14 dpantenna l=0.78u w=0.78u
X2 iovdd.t26 sg13g2_GateDecode_0.pgate.t3 pad.t17 iovdd.t14 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X3 iovdd.t16 sg13g2_GateDecode_0.pgate.t4 pad.t20 iovdd.t14 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X4 iovss sg13g2_GateDecode_0.ngate.t2 pad.t4 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X5 pad.t12 sg13g2_GateDecode_0.pgate.t5 iovdd.t42 iovdd.t14 sg13_hv_pmos ad=3.9294p pd=7.84u as=3.1302p ps=14.26u w=6.66u l=0.6u
X6 iovdd.t22 sg13g2_GateDecode_0.pgate.t6 pad.t15 iovdd.t14 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X7 pad.t22 sg13g2_GateDecode_0.pgate.t7 iovdd.t28 iovdd.t14 sg13_hv_pmos ad=4.9284p pd=14.8u as=2.1312p ps=7.3u w=6.66u l=0.6u
X8 iovss a_12038_31490# p2c.t0 iovss sg13_lv_nmos ad=0.935p pd=6.18u as=0.935p ps=6.18u w=2.75u l=0.13u
X9 iovdd.t27 sg13g2_GateDecode_0.pgate.t4 pad.t19 iovdd.t14 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X10 iovss pad.t25 dantenna l=1.26u w=27.78u
X11 pad.t2 sg13g2_GateDecode_0.ngate.t3 iovss iovss sg13_hv_nmos ad=3.256p pd=10.28u as=1.408p ps=5.04u w=4.4u l=0.6u
X12 pad.t6 sg13g2_GateDecode_0.ngate.t4 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X13 iovss sg13g2_GateDecode_0.ngate.t5 pad.t5 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X14 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t1 c2p_en.t0 a_4230_33842# iovss sg13_lv_nmos ad=1.4148p pd=8.58u as=0.7467p ps=4.31u w=3.93u l=0.13u
X15 iovss sg13g2_LevelDown_0.sg13g2_SecondaryProtection_0.core dantenna l=3.1u w=0.64u
X16 pad.t11 sg13g2_GateDecode_0.pgate.t5 iovdd.t40 iovdd.t14 sg13_hv_pmos ad=3.9294p pd=7.84u as=3.1302p ps=14.26u w=6.66u l=0.6u
X17 iovdd.t15 sg13g2_GateDecode_0.pgate.t6 pad.t14 iovdd.t14 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X18 iovdd.t24 sg13g2_GateDecode_0.pgate.t8 pad.t18 iovdd.t14 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X19 iovss sg13g2_GateDecode_0.ngate.t6 pad.t23 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X20 pad.t21 sg13g2_GateDecode_0.pgate.t7 iovdd.t25 iovdd.t14 sg13_hv_pmos ad=4.9284p pd=14.8u as=2.1312p ps=7.3u w=6.66u l=0.6u
X21 iovdd.t20 sg13g2_GateDecode_0.pgate.t9 pad.t9 iovdd.t14 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X22 iovss sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq iovss sg13_lv_nmos ad=1.4148p pd=8.58u as=0.7467p ps=4.31u w=3.93u l=0.13u
X23 a_12038_31490# sg13g2_LevelDown_0.sg13g2_SecondaryProtection_0.core vdd.t10 vdd.t0 sg13_hv_pmos ad=1.581p pd=9.98u as=1.581p ps=9.98u w=4.65u l=0.45u
X24 a_3724_30170# sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq iovss iovss sg13_hv_nmos ad=0.646p pd=4.48u as=0.361p ps=2.28u w=1.9u l=0.45u
X25 iovdd a_3724_30170# a_3656_30206# iovdd sg13_hv_pmos ad=57f pd=0.68u as=0.102p ps=1.28u w=0.3u l=0.45u
X26 sg13g2_GateDecode_0.ngate.t1 a_3724_30170# iovdd iovdd sg13_hv_pmos ad=1.326p pd=8.48u as=1.326p ps=8.48u w=3.9u l=0.45u
X27 iovdd.t19 sg13g2_GateDecode_0.pgate.t8 pad.t16 iovdd.t14 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X28 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t0 c2p.t0 vdd.t8 vdd.t2 sg13_lv_pmos ad=0.8379p pd=4.79u as=1.4994p ps=9.5u w=4.41u l=0.13u
X29 pad.t20 sg13g2_GateDecode_0.pgate.t10 iovdd.t23 iovdd.t14 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X30 pad.t0 sg13g2_GateDecode_0.ngate.t7 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X31 iovss sg13g2_GateDecode_0.ngate.t8 pad.t3 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X32 pad.t5 sg13g2_GateDecode_0.ngate.t9 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X33 a_4426_30170# a_4358_30206# iovdd iovdd sg13_hv_pmos ad=0.102p pd=1.28u as=57f ps=0.68u w=0.3u l=0.45u
X34 iovdd.t18 sg13g2_GateDecode_0.pgate.t9 pad.t7 iovdd.t14 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X35 a_3750_34876# c2p.t1 vdd.t7 vdd.t6 sg13_lv_pmos ad=0.8379p pd=4.79u as=1.4994p ps=9.5u w=4.41u l=0.13u
X36 pad.t19 sg13g2_GateDecode_0.pgate.t10 iovdd.t17 iovdd.t14 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X37 pad.t8 sg13g2_GateDecode_0.pgate.t11 iovdd.t16 iovdd.t14 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X38 pad.t4 sg13g2_GateDecode_0.ngate.t10 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=2.068p ps=9.74u w=4.4u l=0.6u
X39 pad.t1 sg13g2_GateDecode_0.ngate.t11 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X40 sg13g2_GateDecode_0.ngate.t0 a_3724_30170# iovss iovss sg13_hv_nmos ad=0.646p pd=4.48u as=0.646p ps=4.48u w=1.9u l=0.45u
X41 pad.t18 sg13g2_GateDecode_0.pgate.t12 iovdd.t21 iovdd.t14 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X42 iovdd.t28 sg13g2_GateDecode_0.pgate.t13 pad.t13 iovdd.t14 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X43 vdd.t1 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t2 a_4358_31526# vdd.t0 sg13_lv_pmos ad=1.615p pd=10.18u as=1.615p ps=10.18u w=4.75u l=0.13u
X44 iovss sg13g2_GateDecode_0.ngate.t12 dantenna l=0.78u w=0.78u
X45 iovss a_4358_31526# a_4358_30206# iovss sg13_hv_nmos ad=0.361p pd=2.28u as=0.646p ps=4.48u w=1.9u l=0.45u
X46 pad.t26 iovdd.t0 dpantenna l=1.26u w=27.78u
X47 sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq c2p_en.t1 iovss iovss sg13_lv_nmos ad=1.3362p pd=8.54u as=1.3362p ps=8.54u w=3.93u l=0.13u
X48 iovss sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t2 a_4358_31526# iovss sg13_lv_nmos ad=0.935p pd=6.18u as=0.935p ps=6.18u w=2.75u l=0.13u
X49 pad.t17 sg13g2_GateDecode_0.pgate.t11 iovdd.t27 iovdd.t14 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X50 pad.t16 sg13g2_GateDecode_0.pgate.t12 iovdd.t26 iovdd.t14 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X51 iovss sg13g2_GateDecode_0.ngate.t13 pad.t0 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X52 iovdd.t25 sg13g2_GateDecode_0.pgate.t13 pad.t10 iovdd.t14 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X53 pad.t15 sg13g2_GateDecode_0.pgate.t14 iovdd.t24 iovdd.t14 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X54 vdd.t3 c2p_en.t0 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t0 vdd.t2 sg13_lv_pmos ad=1.5876p pd=9.54u as=0.8379p ps=4.79u w=4.41u l=0.13u
X55 sg13g2_LevelDown_0.sg13g2_SecondaryProtection_0.core pad.t24 iovss rppd l=2u w=1u
X56 iovss sg13g2_GateDecode_0.ngate.t14 pad.t6 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X57 sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq a_3750_34876# vdd.t6 sg13_lv_pmos ad=1.5876p pd=9.54u as=0.8379p ps=4.79u w=4.41u l=0.13u
X58 a_3724_30170# a_3656_30206# iovdd iovdd sg13_hv_pmos ad=0.102p pd=1.28u as=57f ps=0.68u w=0.3u l=0.45u
X59 iovss sg13g2_GateDecode_0.ngate.t15 pad.t1 iovss sg13_hv_nmos ad=1.408p pd=5.04u as=2.596p ps=5.58u w=4.4u l=0.6u
X60 pad.t14 sg13g2_GateDecode_0.pgate.t14 iovdd.t19 iovdd.t14 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X61 pad.t13 sg13g2_GateDecode_0.pgate.t15 iovdd.t20 iovdd.t14 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X62 pad.t27 iovdd.t0 dpantenna l=1.26u w=27.78u
X63 iovdd.t23 sg13g2_GateDecode_0.pgate.t16 pad.t12 iovdd.t14 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X64 sg13g2_GateDecode_0.pgate.t1 a_4426_30170# iovdd iovdd sg13_hv_pmos ad=1.326p pd=8.48u as=1.326p ps=8.48u w=3.9u l=0.45u
X65 pad.t3 sg13g2_GateDecode_0.ngate.t16 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X66 vdd.t9 sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq a_3656_31526# vdd.t0 sg13_lv_pmos ad=1.615p pd=10.18u as=1.615p ps=10.18u w=4.75u l=0.13u
X67 iovss pad.t28 dantenna l=1.26u w=27.78u
X68 a_4230_33842# c2p.t0 iovss iovss sg13_lv_nmos ad=0.7467p pd=4.31u as=1.3362p ps=8.54u w=3.93u l=0.13u
X69 iovss a_3656_31526# a_3656_30206# iovss sg13_hv_nmos ad=0.361p pd=2.28u as=0.646p ps=4.48u w=1.9u l=0.45u
X70 sg13g2_LevelDown_0.sg13g2_SecondaryProtection_0.core iovdd dpantenna l=0.64u w=4.98u
X71 iovdd.t17 sg13g2_GateDecode_0.pgate.t16 pad.t11 iovdd.t14 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X72 pad.t10 sg13g2_GateDecode_0.pgate.t15 iovdd.t18 iovdd.t14 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X73 pad.t9 sg13g2_GateDecode_0.pgate.t17 iovdd.t22 iovdd.t14 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X74 iovdd.t21 sg13g2_GateDecode_0.pgate.t3 pad.t8 iovdd.t14 sg13_hv_pmos ad=2.1312p pd=7.3u as=3.9294p ps=7.84u w=6.66u l=0.6u
X75 iovss sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq a_3656_31526# iovss sg13_lv_nmos ad=0.935p pd=6.18u as=0.935p ps=6.18u w=2.75u l=0.13u
X76 a_4426_30170# sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t3 iovss iovss sg13_hv_nmos ad=0.646p pd=4.48u as=0.361p ps=2.28u w=1.9u l=0.45u
X77 iovdd a_4426_30170# a_4358_30206# iovdd sg13_hv_pmos ad=57f pd=0.68u as=0.102p ps=1.28u w=0.3u l=0.45u
X78 pad.t23 sg13g2_GateDecode_0.ngate.t17 iovss iovss sg13_hv_nmos ad=2.596p pd=5.58u as=1.408p ps=5.04u w=4.4u l=0.6u
X79 sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq c2p.t1 iovss iovss sg13_lv_nmos ad=0.7467p pd=4.31u as=1.3362p ps=8.54u w=3.93u l=0.13u
X80 pad.t7 sg13g2_GateDecode_0.pgate.t17 iovdd.t15 iovdd.t14 sg13_hv_pmos ad=3.9294p pd=7.84u as=2.1312p ps=7.3u w=6.66u l=0.6u
X81 sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq c2p_en.t1 vdd.t5 vdd.t4 sg13_lv_pmos ad=1.4994p pd=9.5u as=1.4994p ps=9.5u w=4.41u l=0.13u
X82 a_12038_31490# sg13g2_LevelDown_0.sg13g2_SecondaryProtection_0.core iovss iovss sg13_hv_nmos ad=0.901p pd=5.98u as=0.901p ps=5.98u w=2.65u l=0.45u
X83 sg13g2_GateDecode_0.pgate.t0 a_4426_30170# iovss iovss sg13_hv_nmos ad=0.646p pd=4.48u as=0.646p ps=4.48u w=1.9u l=0.45u
R0 p2c.n3 p2c 9.10188
R1 p2c.n3 p2c.n2 5.37153
R2 p2c p2c.n3 3.8549
R3 p2c.n0 p2c.t0 1.90938
R4 p2c.n1 p2c.t1 1.76324
R5 p2c.n1 p2c.n0 1.52928
R6 p2c.n2 p2c 1.27498
R7 p2c.n0 p2c 0.673576
R8 p2c.n2 p2c.n1 0.441789
R9 vdd.n39 vdd.n38 23.1683
R10 vdd.n30 vdd.t5 17.0005
R11 vdd.n32 vdd.t3 17.0005
R12 vdd.n34 vdd.t8 17.0005
R13 vdd.n27 vdd.t7 17.0005
R14 vdd.n30 vdd.t4 11.3504
R15 vdd.n37 vdd.t6 11.3229
R16 vdd.n19 vdd.n15 8.45671
R17 vdd.n25 vdd.n15 8.45671
R18 vdd.n22 vdd.n15 8.45671
R19 vdd.n33 vdd.n28 5.65625
R20 vdd.n31 vdd.n28 5.65625
R21 vdd.n36 vdd.n35 5.64342
R22 vdd.n26 vdd.n15 5.58952
R23 vdd.n14 vdd.n13 3.57795
R24 vdd.n41 vdd.n40 3.42019
R25 vdd.n29 vdd.n28 2.83433
R26 vdd.n24 vdd.t9 2.67724
R27 vdd.n21 vdd.t1 2.67724
R28 vdd.n42 vdd.n13 2.5353
R29 vdd.n23 vdd.n15 2.23747
R30 vdd.n20 vdd 2.0602
R31 vdd.n40 vdd.n39 1.94181
R32 vdd.n21 vdd.n20 1.88114
R33 vdd.n16 vdd.n13 1.78381
R34 vdd.n104 vdd.n103 1.50539
R35 vdd.n1 vdd.n0 1.5005
R36 vdd.n99 vdd.n98 1.5005
R37 vdd.n97 vdd.n96 1.5005
R38 vdd.n5 vdd.n4 1.5005
R39 vdd.n91 vdd.n90 1.5005
R40 vdd.n89 vdd.n88 1.5005
R41 vdd.n9 vdd.n8 1.5005
R42 vdd.n83 vdd.n82 1.5005
R43 vdd.n81 vdd.n80 1.5005
R44 vdd.n43 vdd.n12 1.5005
R45 vdd.n75 vdd.n74 1.5005
R46 vdd.n73 vdd.n72 1.5005
R47 vdd.n47 vdd.n46 1.5005
R48 vdd.n67 vdd.n66 1.5005
R49 vdd.n65 vdd.n64 1.5005
R50 vdd.n51 vdd.n50 1.5005
R51 vdd.n59 vdd.n58 1.5005
R52 vdd.n57 vdd.n56 1.5005
R53 vdd.n18 vdd.n16 1.39095
R54 vdd.n17 vdd.t10 1.31928
R55 vdd.n17 vdd.t11 1.21415
R56 vdd.n18 vdd 0.883119
R57 vdd.n23 vdd 0.719451
R58 vdd.n105 vdd 0.6957
R59 vdd.n24 vdd.n23 0.67542
R60 vdd.n103 vdd.n102 0.314786
R61 vdd.n101 vdd.n100 0.314786
R62 vdd.n3 vdd.n2 0.314786
R63 vdd.n95 vdd.n94 0.314786
R64 vdd.n93 vdd.n92 0.314786
R65 vdd.n7 vdd.n6 0.314786
R66 vdd.n87 vdd.n86 0.314786
R67 vdd.n85 vdd.n84 0.314786
R68 vdd.n11 vdd.n10 0.314786
R69 vdd.n79 vdd.n78 0.314786
R70 vdd.n77 vdd.n76 0.314786
R71 vdd.n45 vdd.n44 0.314786
R72 vdd.n71 vdd.n70 0.314786
R73 vdd.n69 vdd.n68 0.314786
R74 vdd.n49 vdd.n48 0.314786
R75 vdd.n63 vdd.n62 0.314786
R76 vdd.n61 vdd.n60 0.314786
R77 vdd.n53 vdd.n52 0.314786
R78 vdd vdd.n22 0.296488
R79 vdd vdd.n25 0.296488
R80 vdd.n39 vdd.n26 0.287915
R81 vdd.n26 vdd 0.264001
R82 vdd vdd.n19 0.249346
R83 vdd vdd.n17 0.233823
R84 vdd.n54 vdd 0.217715
R85 vdd.n55 vdd.n54 0.146103
R86 vdd.n19 vdd.n18 0.110536
R87 vdd.n22 vdd.n21 0.105298
R88 vdd.n25 vdd.n24 0.105298
R89 vdd.n81 vdd.n42 0.0983261
R90 vdd.n35 vdd 0.0934694
R91 vdd.n42 vdd.n41 0.0897467
R92 vdd.n35 vdd.n27 0.0756715
R93 vdd.n14 vdd.t0 0.0745867
R94 vdd.n31 vdd 0.0540006
R95 vdd.n33 vdd.n32 0.0475075
R96 vdd.n37 vdd 0.0474603
R97 vdd.n38 vdd.n37 0.0360492
R98 vdd.n56 vdd.n55 0.0354467
R99 vdd.n34 vdd.n33 0.0348561
R100 vdd.n32 vdd.n31 0.0333284
R101 vdd.n55 vdd.n52 0.0314255
R102 vdd vdd.n30 0.0199792
R103 vdd vdd.n34 0.0199792
R104 vdd.n27 vdd 0.0199792
R105 vdd.n40 vdd.n15 0.0167109
R106 vdd.n16 vdd.n15 0.0155555
R107 vdd.n18 vdd 0.01205
R108 vdd.n38 vdd 0.0115764
R109 vdd.n58 vdd.n57 0.00921287
R110 vdd.n58 vdd.n50 0.00921287
R111 vdd.n65 vdd.n50 0.00921287
R112 vdd.n66 vdd.n65 0.00921287
R113 vdd.n66 vdd.n46 0.00921287
R114 vdd.n73 vdd.n46 0.00921287
R115 vdd.n74 vdd.n73 0.00921287
R116 vdd.n74 vdd.n12 0.00921287
R117 vdd.n81 vdd.n12 0.00921287
R118 vdd.n82 vdd.n81 0.00921287
R119 vdd.n82 vdd.n8 0.00921287
R120 vdd.n89 vdd.n8 0.00921287
R121 vdd.n90 vdd.n89 0.00921287
R122 vdd.n90 vdd.n4 0.00921287
R123 vdd.n97 vdd.n4 0.00921287
R124 vdd.n98 vdd.n97 0.00921287
R125 vdd.n98 vdd.n0 0.00921287
R126 vdd.n104 vdd.n0 0.00921287
R127 vdd.n41 vdd 0.00903111
R128 vdd.n56 vdd.n53 0.00538889
R129 vdd.n59 vdd.n53 0.00538889
R130 vdd.n60 vdd.n59 0.00538889
R131 vdd.n60 vdd.n51 0.00538889
R132 vdd.n63 vdd.n51 0.00538889
R133 vdd.n64 vdd.n63 0.00538889
R134 vdd.n64 vdd.n49 0.00538889
R135 vdd.n67 vdd.n49 0.00538889
R136 vdd.n68 vdd.n67 0.00538889
R137 vdd.n68 vdd.n47 0.00538889
R138 vdd.n71 vdd.n47 0.00538889
R139 vdd.n72 vdd.n71 0.00538889
R140 vdd.n72 vdd.n45 0.00538889
R141 vdd.n75 vdd.n45 0.00538889
R142 vdd.n76 vdd.n75 0.00538889
R143 vdd.n76 vdd.n43 0.00538889
R144 vdd.n79 vdd.n43 0.00538889
R145 vdd.n80 vdd.n79 0.00538889
R146 vdd.n80 vdd.n11 0.00538889
R147 vdd.n83 vdd.n11 0.00538889
R148 vdd.n84 vdd.n83 0.00538889
R149 vdd.n84 vdd.n9 0.00538889
R150 vdd.n87 vdd.n9 0.00538889
R151 vdd.n88 vdd.n87 0.00538889
R152 vdd.n88 vdd.n7 0.00538889
R153 vdd.n91 vdd.n7 0.00538889
R154 vdd.n92 vdd.n91 0.00538889
R155 vdd.n92 vdd.n5 0.00538889
R156 vdd.n95 vdd.n5 0.00538889
R157 vdd.n96 vdd.n95 0.00538889
R158 vdd.n96 vdd.n3 0.00538889
R159 vdd.n99 vdd.n3 0.00538889
R160 vdd.n100 vdd.n99 0.00538889
R161 vdd.n100 vdd.n1 0.00538889
R162 vdd.n103 vdd.n1 0.00538889
R163 vdd.n57 vdd.n54 0.00485644
R164 vdd.n105 vdd.n104 0.00485644
R165 vdd vdd.n105 0.00485644
R166 vdd.n102 vdd 0.0035
R167 vdd.n61 vdd.n52 0.0025
R168 vdd.n62 vdd.n61 0.0025
R169 vdd.n62 vdd.n48 0.0025
R170 vdd.n69 vdd.n48 0.0025
R171 vdd.n70 vdd.n69 0.0025
R172 vdd.n70 vdd.n44 0.0025
R173 vdd.n77 vdd.n44 0.0025
R174 vdd.n78 vdd.n77 0.0025
R175 vdd.n78 vdd.n10 0.0025
R176 vdd.n85 vdd.n10 0.0025
R177 vdd.n86 vdd.n85 0.0025
R178 vdd.n86 vdd.n6 0.0025
R179 vdd.n93 vdd.n6 0.0025
R180 vdd.n94 vdd.n93 0.0025
R181 vdd.n94 vdd.n2 0.0025
R182 vdd.n101 vdd.n2 0.0025
R183 vdd.n102 vdd.n101 0.0025
R184 vdd.n20 vdd.n15 0.00245557
R185 vdd.n15 vdd.n14 0.00100649
R186 vdd.n29 vdd.t2 0.001
R187 vdd.t6 vdd.n36 0.001
R188 vdd.t4 vdd.n29 0.001
R189 vdd.n36 vdd.t2 0.001
R190 sg13g2_GateDecode_0.sg13g2_LevelUp_1.o sg13g2_GateDecode_0.pgate.n18 32.6396
R191 sg13g2_GateDecode_0.pgate.n17 sg13g2_GateDecode_0.pgate.n15 9.58949
R192 sg13g2_GateDecode_0.pgate.n16 sg13g2_GateDecode_0.pgate.n1 9.00605
R193 sg13g2_GateDecode_0.pgate.n18 sg13g2_GateDecode_0.pgate.n17 9.0005
R194 sg13g2_GateDecode_0.pgate.n2 sg13g2_GateDecode_0.pgate.t7 7.94005
R195 sg13g2_GateDecode_0.pgate.n15 sg13g2_GateDecode_0.pgate.t5 7.08755
R196 sg13g2_GateDecode_0.pgate.n2 sg13g2_GateDecode_0.pgate.t13 7.08755
R197 sg13g2_GateDecode_0.pgate.n3 sg13g2_GateDecode_0.pgate.t15 7.08755
R198 sg13g2_GateDecode_0.pgate.n4 sg13g2_GateDecode_0.pgate.t9 7.08755
R199 sg13g2_GateDecode_0.pgate.n5 sg13g2_GateDecode_0.pgate.t17 7.08755
R200 sg13g2_GateDecode_0.pgate.n6 sg13g2_GateDecode_0.pgate.t6 7.08755
R201 sg13g2_GateDecode_0.pgate.n7 sg13g2_GateDecode_0.pgate.t14 7.08755
R202 sg13g2_GateDecode_0.pgate.n8 sg13g2_GateDecode_0.pgate.t8 7.08755
R203 sg13g2_GateDecode_0.pgate.n9 sg13g2_GateDecode_0.pgate.t12 7.08755
R204 sg13g2_GateDecode_0.pgate.n10 sg13g2_GateDecode_0.pgate.t3 7.08755
R205 sg13g2_GateDecode_0.pgate.n11 sg13g2_GateDecode_0.pgate.t11 7.08755
R206 sg13g2_GateDecode_0.pgate.n12 sg13g2_GateDecode_0.pgate.t4 7.08755
R207 sg13g2_GateDecode_0.pgate.n13 sg13g2_GateDecode_0.pgate.t10 7.08755
R208 sg13g2_GateDecode_0.pgate.n14 sg13g2_GateDecode_0.pgate.t16 7.08755
R209 sg13g2_GateDecode_0.pgate.n0 sg13g2_GateDecode_0.pgate.t0 4.59834
R210 sg13g2_GateDecode_0.pgate.n16 sg13g2_GateDecode_0.pgate.t2 4.2615
R211 sg13g2_GateDecode_0.pgate.n0 sg13g2_GateDecode_0.pgate.t1 2.00385
R212 sg13g2_GateDecode_0.sg13g2_LevelUp_1.o sg13g2_GateDecode_0.pgate.n0 1.98894
R213 sg13g2_GateDecode_0.pgate.n3 sg13g2_GateDecode_0.pgate.n2 1.22425
R214 sg13g2_GateDecode_0.pgate.n5 sg13g2_GateDecode_0.pgate.n4 1.22425
R215 sg13g2_GateDecode_0.pgate.n7 sg13g2_GateDecode_0.pgate.n6 1.22425
R216 sg13g2_GateDecode_0.pgate.n9 sg13g2_GateDecode_0.pgate.n8 1.22425
R217 sg13g2_GateDecode_0.pgate.n11 sg13g2_GateDecode_0.pgate.n10 1.22425
R218 sg13g2_GateDecode_0.pgate.n13 sg13g2_GateDecode_0.pgate.n12 1.22425
R219 sg13g2_GateDecode_0.pgate.n15 sg13g2_GateDecode_0.pgate.n14 1.22425
R220 sg13g2_GateDecode_0.pgate.n4 sg13g2_GateDecode_0.pgate.n3 0.853
R221 sg13g2_GateDecode_0.pgate.n6 sg13g2_GateDecode_0.pgate.n5 0.853
R222 sg13g2_GateDecode_0.pgate.n8 sg13g2_GateDecode_0.pgate.n7 0.853
R223 sg13g2_GateDecode_0.pgate.n10 sg13g2_GateDecode_0.pgate.n9 0.853
R224 sg13g2_GateDecode_0.pgate.n12 sg13g2_GateDecode_0.pgate.n11 0.853
R225 sg13g2_GateDecode_0.pgate.n14 sg13g2_GateDecode_0.pgate.n13 0.853
R226 sg13g2_GateDecode_0.pgate.n18 sg13g2_GateDecode_0.pgate.n1 0.2117
R227 sg13g2_GateDecode_0.pgate.n17 sg13g2_GateDecode_0.pgate.n16 0.201404
R228 sg13g2_GateDecode_0.pgate.n1 sg13g2_Clamp_P15N15D_0.gate 0.0841
R229 iovdd.n305 iovdd.n304 10.8089
R230 iovdd.n299 iovdd.n298 10.8089
R231 iovdd.n268 iovdd.n267 10.8089
R232 iovdd.n244 iovdd.n243 10.8089
R233 iovdd.n241 iovdd.n240 10.8089
R234 iovdd.n271 iovdd.n270 10.8089
R235 iovdd.n302 iovdd.n120 10.8089
R236 iovdd.n264 iovdd.n263 10.8089
R237 iovdd.n277 iovdd.n276 9.0005
R238 iovdd.n445 iovdd.n444 9.0005
R239 iovdd.n442 iovdd.n441 9.0005
R240 iovdd.n427 iovdd.n426 9.0005
R241 iovdd.n236 iovdd.n30 9.0005
R242 iovdd.n468 iovdd.n467 9.0005
R243 iovdd.n424 iovdd.n423 9.0005
R244 iovdd.n465 iovdd.n464 9.0005
R245 iovdd.n500 iovdd.n31 5.66717
R246 iovdd.n501 iovdd.n500 5.66717
R247 iovdd.n457 iovdd.n456 5.66717
R248 iovdd.n456 iovdd.n455 5.66717
R249 iovdd.n437 iovdd.n111 5.66717
R250 iovdd.n438 iovdd.n437 5.66717
R251 iovdd.n419 iovdd.n407 5.66717
R252 iovdd.n420 iovdd.n419 5.66717
R253 iovdd.n415 iovdd.n414 5.66717
R254 iovdd.n414 iovdd.n413 5.66717
R255 iovdd.n430 iovdd.n428 4.9805
R256 iovdd.n104 iovdd.n102 4.9805
R257 iovdd.n448 iovdd.n446 4.9805
R258 iovdd.n471 iovdd.n469 4.9805
R259 iovdd.n506 iovdd.n505 4.9805
R260 iovdd.n274 iovdd.n272 4.9805
R261 iovdd.n80 iovdd.n78 4.9805
R262 iovdd.n509 iovdd.n21 4.28068
R263 iovdd.n511 iovdd.n18 4.2505
R264 iovdd.n398 iovdd.n396 3.0005
R265 iovdd.n400 iovdd.n395 3.0005
R266 iovdd.n430 iovdd.n429 3.0005
R267 iovdd.n104 iovdd.n103 3.0005
R268 iovdd.n448 iovdd.n447 3.0005
R269 iovdd.n274 iovdd.n273 3.0005
R270 iovdd.n471 iovdd.n470 3.0005
R271 iovdd.n505 iovdd.n504 3.0005
R272 iovdd.n422 iovdd.n421 3.0005
R273 iovdd.n432 iovdd.n431 3.0005
R274 iovdd.n440 iovdd.n439 3.0005
R275 iovdd.n450 iovdd.n449 3.0005
R276 iovdd.n275 iovdd.n91 3.0005
R277 iovdd.n473 iovdd.n472 3.0005
R278 iovdd.n503 iovdd.n502 3.0005
R279 iovdd.n463 iovdd.n462 3.0005
R280 iovdd.n80 iovdd.n79 3.0005
R281 iovdd.t0 iovdd.n498 2.83433
R282 iovdd.t0 iovdd.n483 2.83433
R283 iovdd.t0 iovdd.n482 2.83433
R284 iovdd.t0 iovdd.n481 2.83433
R285 iovdd.t0 iovdd.n480 2.83433
R286 iovdd.t0 iovdd.n479 2.83433
R287 iovdd.t0 iovdd.n33 2.83433
R288 iovdd.n499 iovdd.t0 2.83433
R289 iovdd.t0 iovdd.n478 2.83433
R290 iovdd.t0 iovdd.n68 2.83433
R291 iovdd.t0 iovdd.n67 2.83433
R292 iovdd.t0 iovdd.n66 2.83433
R293 iovdd.t0 iovdd.n65 2.83433
R294 iovdd.t0 iovdd.n64 2.83433
R295 iovdd.t0 iovdd.n63 2.83433
R296 iovdd.t0 iovdd.n62 2.83433
R297 iovdd.t0 iovdd.n61 2.83433
R298 iovdd.t0 iovdd.n60 2.83433
R299 iovdd.t0 iovdd.n59 2.83433
R300 iovdd.t0 iovdd.n58 2.83433
R301 iovdd.t0 iovdd.n57 2.83433
R302 iovdd.t0 iovdd.n56 2.83433
R303 iovdd.t0 iovdd.n55 2.83433
R304 iovdd.t0 iovdd.n54 2.83433
R305 iovdd.t0 iovdd.n53 2.83433
R306 iovdd.t0 iovdd.n52 2.83433
R307 iovdd.t0 iovdd.n51 2.83433
R308 iovdd.t0 iovdd.n50 2.83433
R309 iovdd.t0 iovdd.n49 2.83433
R310 iovdd.t0 iovdd.n48 2.83433
R311 iovdd.t0 iovdd.n47 2.83433
R312 iovdd.t0 iovdd.n46 2.83433
R313 iovdd.t0 iovdd.n45 2.83433
R314 iovdd.t0 iovdd.n44 2.83433
R315 iovdd.t0 iovdd.n43 2.83433
R316 iovdd.t0 iovdd.n42 2.83433
R317 iovdd.t0 iovdd.n41 2.83433
R318 iovdd.t0 iovdd.n40 2.83433
R319 iovdd.t0 iovdd.n39 2.83433
R320 iovdd.t0 iovdd.n38 2.83433
R321 iovdd.t0 iovdd.n37 2.83433
R322 iovdd.t0 iovdd.n36 2.83433
R323 iovdd.n497 iovdd.n496 2.82693
R324 iovdd.n495 iovdd.n484 2.82693
R325 iovdd.n494 iovdd.n485 2.82693
R326 iovdd.n493 iovdd.n486 2.82693
R327 iovdd.n492 iovdd.n487 2.82693
R328 iovdd.n491 iovdd.n488 2.82693
R329 iovdd.n490 iovdd.n489 2.82693
R330 iovdd.n34 iovdd.n32 2.82693
R331 iovdd.n477 iovdd.n476 2.82693
R332 iovdd.n475 iovdd.n69 2.82693
R333 iovdd.n474 iovdd.n70 2.82693
R334 iovdd.n72 iovdd.n71 2.82693
R335 iovdd.n82 iovdd.n81 2.82693
R336 iovdd.n84 iovdd.n83 2.82693
R337 iovdd.n86 iovdd.n85 2.82693
R338 iovdd.n461 iovdd.n87 2.82693
R339 iovdd.n460 iovdd.n88 2.82693
R340 iovdd.n459 iovdd.n89 2.82693
R341 iovdd.n458 iovdd.n90 2.82693
R342 iovdd.n454 iovdd.n92 2.82693
R343 iovdd.n453 iovdd.n93 2.82693
R344 iovdd.n452 iovdd.n94 2.82693
R345 iovdd.n451 iovdd.n95 2.82693
R346 iovdd.n97 iovdd.n96 2.82693
R347 iovdd.n106 iovdd.n105 2.82693
R348 iovdd.n108 iovdd.n107 2.82693
R349 iovdd.n110 iovdd.n109 2.82693
R350 iovdd.n436 iovdd.n112 2.82693
R351 iovdd.n435 iovdd.n113 2.82693
R352 iovdd.n434 iovdd.n114 2.82693
R353 iovdd.n433 iovdd.n115 2.82693
R354 iovdd.n117 iovdd.n116 2.82693
R355 iovdd.n402 iovdd.n401 2.82693
R356 iovdd.n404 iovdd.n403 2.82693
R357 iovdd.n406 iovdd.n405 2.82693
R358 iovdd.n418 iovdd.n408 2.82693
R359 iovdd.n417 iovdd.n409 2.82693
R360 iovdd.n416 iovdd.n410 2.82693
R361 iovdd.n511 iovdd.n2 2.41731
R362 iovdd.n512 iovdd.n511 2.1192
R363 iovdd.n511 iovdd.n15 2.11861
R364 iovdd.n100 iovdd.n75 1.98828
R365 iovdd.n300 iovdd.n75 1.98792
R366 iovdd.n431 iovdd.n430 1.9805
R367 iovdd.n440 iovdd.n104 1.9805
R368 iovdd.n449 iovdd.n448 1.9805
R369 iovdd.n472 iovdd.n471 1.9805
R370 iovdd.n505 iovdd.n503 1.9805
R371 iovdd.n275 iovdd.n274 1.9805
R372 iovdd.n463 iovdd.n80 1.9805
R373 iovdd.t0 iovdd.n35 1.89
R374 iovdd.n431 iovdd.n427 1.8749
R375 iovdd.n441 iovdd.n440 1.8749
R376 iovdd.n449 iovdd.n445 1.8749
R377 iovdd.n472 iovdd.n468 1.8749
R378 iovdd.n503 iovdd.n30 1.8749
R379 iovdd.n277 iovdd.n275 1.8749
R380 iovdd.n464 iovdd.n463 1.8749
R381 iovdd.n427 iovdd.n118 1.8089
R382 iovdd.n441 iovdd.n101 1.8089
R383 iovdd.n445 iovdd.n98 1.8089
R384 iovdd.n468 iovdd.n73 1.8089
R385 iovdd.n238 iovdd.n30 1.8089
R386 iovdd.n278 iovdd.n277 1.8089
R387 iovdd.n423 iovdd.n393 1.8089
R388 iovdd.n464 iovdd.n77 1.8089
R389 iovdd.n263 iovdd.t15 1.76518
R390 iovdd.n77 iovdd.t22 1.76518
R391 iovdd.n271 iovdd.t19 1.76518
R392 iovdd.n278 iovdd.t24 1.76518
R393 iovdd.n305 iovdd.t17 1.76518
R394 iovdd.n118 iovdd.t23 1.76518
R395 iovdd.n298 iovdd.t27 1.76518
R396 iovdd.n101 iovdd.t16 1.76518
R397 iovdd.n267 iovdd.t26 1.76518
R398 iovdd.n98 iovdd.t21 1.76518
R399 iovdd.n244 iovdd.t18 1.76518
R400 iovdd.n73 iovdd.t20 1.76518
R401 iovdd.n240 iovdd.t25 1.76518
R402 iovdd.n238 iovdd.t28 1.76518
R403 iovdd.n120 iovdd.t40 1.76484
R404 iovdd.n393 iovdd.t42 1.76484
R405 iovdd.n425 iovdd.n75 1.73634
R406 iovdd.n99 iovdd.n75 1.73634
R407 iovdd.n466 iovdd.n75 1.73634
R408 iovdd.n443 iovdd.n75 1.73611
R409 iovdd.n76 iovdd.n75 1.73611
R410 iovdd.n75 iovdd.n74 1.73611
R411 iovdd.n133 iovdd.n75 1.73611
R412 iovdd.n265 iovdd.n75 1.73611
R413 iovdd.n242 iovdd.n75 1.73611
R414 iovdd.n303 iovdd.n75 1.73595
R415 iovdd.n269 iovdd.n75 1.73595
R416 iovdd.n144 iovdd.n75 1.73595
R417 iovdd.t0 iovdd.n1 1.70106
R418 iovdd.n412 iovdd.n411 1.68243
R419 iovdd.n423 iovdd.n422 1.60815
R420 iovdd.n306 iovdd.n305 1.5625
R421 iovdd.n306 iovdd.n118 1.5625
R422 iovdd.n298 iovdd.n297 1.5625
R423 iovdd.n297 iovdd.n101 1.5625
R424 iovdd.n267 iovdd.n266 1.5625
R425 iovdd.n266 iovdd.n98 1.5625
R426 iovdd.n245 iovdd.n244 1.5625
R427 iovdd.n245 iovdd.n73 1.5625
R428 iovdd.n240 iovdd.n239 1.5625
R429 iovdd.n239 iovdd.n238 1.5625
R430 iovdd.n279 iovdd.n271 1.5625
R431 iovdd.n279 iovdd.n278 1.5625
R432 iovdd.n392 iovdd.n120 1.5625
R433 iovdd.n393 iovdd.n392 1.5625
R434 iovdd.n263 iovdd.n262 1.5625
R435 iovdd.n262 iovdd.n77 1.5625
R436 iovdd iovdd.n119 1.43219
R437 iovdd.n241 iovdd.n237 1.42534
R438 iovdd.n237 iovdd.n236 1.42433
R439 iovdd.n301 iovdd 1.39634
R440 iovdd.n424 iovdd.n119 1.33976
R441 iovdd.n302 iovdd.n301 1.33311
R442 iovdd.n511 iovdd.n14 1.28534
R443 iovdd.n511 iovdd.n20 1.28534
R444 iovdd.n355 iovdd.n351 0.826084
R445 iovdd.n188 iovdd.n181 0.826084
R446 iovdd.n358 iovdd.n350 0.818682
R447 iovdd.n349 iovdd.n342 0.818682
R448 iovdd.n365 iovdd.n341 0.818682
R449 iovdd.n366 iovdd.n340 0.818682
R450 iovdd.n339 iovdd.n332 0.818682
R451 iovdd.n373 iovdd.n331 0.818682
R452 iovdd.n374 iovdd.n330 0.818682
R453 iovdd.n329 iovdd.n322 0.818682
R454 iovdd.n381 iovdd.n321 0.818682
R455 iovdd.n382 iovdd.n320 0.818682
R456 iovdd.n124 iovdd.n122 0.818682
R457 iovdd.n390 iovdd.n389 0.818682
R458 iovdd.n123 iovdd.n121 0.818682
R459 iovdd.n309 iovdd.n308 0.818682
R460 iovdd.n132 iovdd.n131 0.818682
R461 iovdd.n295 iovdd.n294 0.818682
R462 iovdd.n281 iovdd.n135 0.818682
R463 iovdd.n283 iovdd.n282 0.818682
R464 iovdd.n143 iovdd.n142 0.818682
R465 iovdd.n260 iovdd.n259 0.818682
R466 iovdd.n146 iovdd.n145 0.818682
R467 iovdd.n248 iovdd.n247 0.818682
R468 iovdd.n234 iovdd.n153 0.818682
R469 iovdd.n233 iovdd.n232 0.818682
R470 iovdd.n155 iovdd.n154 0.818682
R471 iovdd.n221 iovdd.n220 0.818682
R472 iovdd.n219 iovdd.n162 0.818682
R473 iovdd.n218 iovdd.n217 0.818682
R474 iovdd.n164 iovdd.n163 0.818682
R475 iovdd.n206 iovdd.n205 0.818682
R476 iovdd.n204 iovdd.n171 0.818682
R477 iovdd.n203 iovdd.n202 0.818682
R478 iovdd.n173 iovdd.n172 0.818682
R479 iovdd.n191 iovdd.n190 0.818682
R480 iovdd.n189 iovdd.n180 0.818682
R481 iovdd.n187 iovdd.n186 0.818682
R482 iovdd.n182 iovdd.n180 0.818682
R483 iovdd.n192 iovdd.n191 0.818682
R484 iovdd.n193 iovdd.n173 0.818682
R485 iovdd.n202 iovdd.n201 0.818682
R486 iovdd.n175 iovdd.n171 0.818682
R487 iovdd.n207 iovdd.n206 0.818682
R488 iovdd.n208 iovdd.n164 0.818682
R489 iovdd.n217 iovdd.n216 0.818682
R490 iovdd.n166 iovdd.n162 0.818682
R491 iovdd.n222 iovdd.n221 0.818682
R492 iovdd.n223 iovdd.n155 0.818682
R493 iovdd.n232 iovdd.n231 0.818682
R494 iovdd.n157 iovdd.n153 0.818682
R495 iovdd.n249 iovdd.n248 0.818682
R496 iovdd.n250 iovdd.n146 0.818682
R497 iovdd.n259 iovdd.n258 0.818682
R498 iovdd.n148 iovdd.n142 0.818682
R499 iovdd.n284 iovdd.n283 0.818682
R500 iovdd.n285 iovdd.n135 0.818682
R501 iovdd.n294 iovdd.n293 0.818682
R502 iovdd.n137 iovdd.n131 0.818682
R503 iovdd.n310 iovdd.n309 0.818682
R504 iovdd.n311 iovdd.n123 0.818682
R505 iovdd.n389 iovdd.n388 0.818682
R506 iovdd.n126 iovdd.n124 0.818682
R507 iovdd.n383 iovdd.n382 0.818682
R508 iovdd.n381 iovdd.n380 0.818682
R509 iovdd.n323 iovdd.n322 0.818682
R510 iovdd.n375 iovdd.n374 0.818682
R511 iovdd.n373 iovdd.n372 0.818682
R512 iovdd.n333 iovdd.n332 0.818682
R513 iovdd.n367 iovdd.n366 0.818682
R514 iovdd.n365 iovdd.n364 0.818682
R515 iovdd.n343 iovdd.n342 0.818682
R516 iovdd.n359 iovdd.n358 0.818682
R517 iovdd.n357 iovdd.n356 0.818682
R518 iovdd.n511 iovdd.n22 0.671789
R519 iovdd.n511 iovdd.n6 0.671602
R520 iovdd.n511 iovdd.n28 0.671602
R521 iovdd.n511 iovdd.n12 0.671423
R522 iovdd.n511 iovdd.n24 0.588672
R523 iovdd.n511 iovdd.n26 0.588672
R524 iovdd.n511 iovdd.n29 0.588672
R525 iovdd.n511 iovdd.n11 0.588437
R526 iovdd.n511 iovdd.n9 0.588437
R527 iovdd.n511 iovdd.n7 0.588437
R528 iovdd.n511 iovdd.n23 0.588437
R529 iovdd.n511 iovdd.n25 0.588437
R530 iovdd.n511 iovdd.n27 0.588437
R531 iovdd.n511 iovdd.n10 0.588281
R532 iovdd.n511 iovdd.n8 0.588281
R533 iovdd.n511 iovdd.n5 0.588281
R534 iovdd.n511 iovdd.n3 0.588266
R535 iovdd.n444 iovdd.n443 0.515695
R536 iovdd.n268 iovdd.n133 0.515695
R537 iovdd.n425 iovdd.n424 0.513735
R538 iovdd.n303 iovdd.n302 0.513312
R539 iovdd.n511 iovdd.n510 0.503491
R540 iovdd.n270 iovdd.n269 0.502871
R541 iovdd.n276 iovdd.n99 0.502476
R542 iovdd.n511 iovdd.n17 0.502128
R543 iovdd.n465 iovdd.n76 0.489812
R544 iovdd.n265 iovdd.n264 0.489812
R545 iovdd.n467 iovdd.n74 0.481088
R546 iovdd.n243 iovdd.n242 0.481088
R547 iovdd.n300 iovdd.n299 0.479418
R548 iovdd.n442 iovdd.n100 0.479034
R549 iovdd.n426 iovdd.n100 0.477001
R550 iovdd.n243 iovdd.n144 0.476989
R551 iovdd.n304 iovdd.n300 0.476595
R552 iovdd.n467 iovdd.n466 0.476594
R553 iovdd.n466 iovdd.n465 0.468441
R554 iovdd.n264 iovdd.n144 0.468018
R555 iovdd.n236 iovdd.n74 0.46393
R556 iovdd.n242 iovdd.n241 0.46393
R557 iovdd.n276 iovdd.n76 0.455206
R558 iovdd.n270 iovdd.n265 0.455206
R559 iovdd.n444 iovdd.n99 0.442559
R560 iovdd.n269 iovdd.n268 0.442135
R561 iovdd.n304 iovdd.n303 0.431695
R562 iovdd.n426 iovdd.n425 0.4313
R563 iovdd.n443 iovdd.n442 0.429323
R564 iovdd.n299 iovdd.n133 0.429323
R565 iovdd.n189 iovdd.n188 0.416993
R566 iovdd.n351 iovdd.n350 0.416993
R567 iovdd.n507 iovdd.n506 0.328683
R568 iovdd.n508 iovdd.n507 0.270343
R569 iovdd.n508 iovdd.n4 0.258522
R570 iovdd.n511 iovdd.n4 0.254672
R571 iovdd.n398 iovdd.n397 0.2505
R572 iovdd.n400 iovdd.n399 0.2505
R573 iovdd.n422 iovdd.n394 0.2505
R574 iovdd.n504 iovdd.n4 0.227256
R575 iovdd.n183 iovdd.n181 0.201704
R576 iovdd.n355 iovdd.n354 0.2005
R577 iovdd.n348 iovdd.n347 0.2005
R578 iovdd.n361 iovdd.n360 0.2005
R579 iovdd.n363 iovdd.n362 0.2005
R580 iovdd.n338 iovdd.n337 0.2005
R581 iovdd.n369 iovdd.n368 0.2005
R582 iovdd.n371 iovdd.n370 0.2005
R583 iovdd.n328 iovdd.n327 0.2005
R584 iovdd.n377 iovdd.n376 0.2005
R585 iovdd.n379 iovdd.n378 0.2005
R586 iovdd.n319 iovdd.n318 0.2005
R587 iovdd.n385 iovdd.n384 0.2005
R588 iovdd.n387 iovdd.n386 0.2005
R589 iovdd.n127 iovdd.n125 0.2005
R590 iovdd.n313 iovdd.n312 0.2005
R591 iovdd.n130 iovdd.n129 0.2005
R592 iovdd.n292 iovdd.n291 0.2005
R593 iovdd.n138 iovdd.n136 0.2005
R594 iovdd.n287 iovdd.n286 0.2005
R595 iovdd.n141 iovdd.n140 0.2005
R596 iovdd.n257 iovdd.n256 0.2005
R597 iovdd.n149 iovdd.n147 0.2005
R598 iovdd.n252 iovdd.n251 0.2005
R599 iovdd.n152 iovdd.n151 0.2005
R600 iovdd.n230 iovdd.n229 0.2005
R601 iovdd.n158 iovdd.n156 0.2005
R602 iovdd.n225 iovdd.n224 0.2005
R603 iovdd.n161 iovdd.n160 0.2005
R604 iovdd.n215 iovdd.n214 0.2005
R605 iovdd.n167 iovdd.n165 0.2005
R606 iovdd.n210 iovdd.n209 0.2005
R607 iovdd.n170 iovdd.n169 0.2005
R608 iovdd.n200 iovdd.n199 0.2005
R609 iovdd.n176 iovdd.n174 0.2005
R610 iovdd.n195 iovdd.n194 0.2005
R611 iovdd.n179 iovdd.n178 0.2005
R612 iovdd.n185 iovdd.n184 0.2005
R613 iovdd.n262 iovdd.n261 0.191989
R614 iovdd.n280 iovdd.n279 0.191989
R615 iovdd.n266 iovdd.n134 0.191989
R616 iovdd.n297 iovdd.n296 0.191989
R617 iovdd.n307 iovdd.n306 0.191989
R618 iovdd.n392 iovdd.n391 0.191989
R619 iovdd.n239 iovdd.n235 0.191989
R620 iovdd.n246 iovdd.n245 0.191989
R621 iovdd.n17 iovdd.n16 0.156542
R622 iovdd.n510 iovdd.n508 0.153056
R623 iovdd.n3 iovdd.n0 0.144604
R624 iovdd.n504 iovdd.n5 0.143944
R625 iovdd.n506 iovdd.n29 0.14355
R626 iovdd.n272 iovdd.n27 0.142174
R627 iovdd.n273 iovdd.n7 0.142174
R628 iovdd.n16 iovdd.n3 0.139796
R629 iovdd.n446 iovdd.n26 0.138974
R630 iovdd.n447 iovdd.n8 0.138556
R631 iovdd.n102 iovdd.n25 0.13519
R632 iovdd.n103 iovdd.n9 0.13519
R633 iovdd.n429 iovdd.n11 0.135097
R634 iovdd.n428 iovdd.n23 0.135097
R635 iovdd.n470 iovdd.n6 0.133441
R636 iovdd.n469 iovdd.n28 0.133441
R637 iovdd.n428 iovdd.n24 0.13199
R638 iovdd.n103 iovdd.n10 0.131722
R639 iovdd.n78 iovdd.n28 0.131626
R640 iovdd.n79 iovdd.n6 0.131626
R641 iovdd.n429 iovdd.n10 0.131572
R642 iovdd.n102 iovdd.n24 0.131328
R643 iovdd.n396 iovdd.n23 0.128206
R644 iovdd.n395 iovdd.n11 0.128206
R645 iovdd.n447 iovdd.n9 0.128113
R646 iovdd.n446 iovdd.n25 0.128113
R647 iovdd.n510 iovdd.n509 0.127471
R648 iovdd.n395 iovdd.n12 0.124896
R649 iovdd.n273 iovdd.n8 0.124738
R650 iovdd.n19 iovdd.n17 0.124655
R651 iovdd.n396 iovdd.n22 0.124514
R652 iovdd.n272 iovdd.n26 0.124344
R653 iovdd.n79 iovdd.n7 0.121129
R654 iovdd.n78 iovdd.n27 0.121129
R655 iovdd.n469 iovdd.n29 0.119767
R656 iovdd.n470 iovdd.n5 0.11935
R657 iovdd.n397 iovdd.n22 0.117846
R658 iovdd.n399 iovdd.n12 0.117444
R659 iovdd.n354 iovdd.n353 0.1105
R660 iovdd.n352 iovdd.n347 0.1105
R661 iovdd.n361 iovdd.n346 0.1105
R662 iovdd.n362 iovdd.n345 0.1105
R663 iovdd.n344 iovdd.n337 0.1105
R664 iovdd.n369 iovdd.n336 0.1105
R665 iovdd.n370 iovdd.n335 0.1105
R666 iovdd.n334 iovdd.n327 0.1105
R667 iovdd.n377 iovdd.n326 0.1105
R668 iovdd.n378 iovdd.n325 0.1105
R669 iovdd.n324 iovdd.n318 0.1105
R670 iovdd.n385 iovdd.n317 0.1105
R671 iovdd.n386 iovdd.n316 0.1105
R672 iovdd.n315 iovdd.n127 0.1105
R673 iovdd.n314 iovdd.n313 0.1105
R674 iovdd.n129 iovdd.n128 0.1105
R675 iovdd.n291 iovdd.n290 0.1105
R676 iovdd.n289 iovdd.n138 0.1105
R677 iovdd.n288 iovdd.n287 0.1105
R678 iovdd.n140 iovdd.n139 0.1105
R679 iovdd.n256 iovdd.n255 0.1105
R680 iovdd.n254 iovdd.n149 0.1105
R681 iovdd.n253 iovdd.n252 0.1105
R682 iovdd.n151 iovdd.n150 0.1105
R683 iovdd.n229 iovdd.n228 0.1105
R684 iovdd.n227 iovdd.n158 0.1105
R685 iovdd.n226 iovdd.n225 0.1105
R686 iovdd.n160 iovdd.n159 0.1105
R687 iovdd.n214 iovdd.n213 0.1105
R688 iovdd.n212 iovdd.n167 0.1105
R689 iovdd.n211 iovdd.n210 0.1105
R690 iovdd.n169 iovdd.n168 0.1105
R691 iovdd.n199 iovdd.n198 0.1105
R692 iovdd.n197 iovdd.n176 0.1105
R693 iovdd.n196 iovdd.n195 0.1105
R694 iovdd.n178 iovdd.n177 0.1105
R695 iovdd.n511 iovdd.n507 0.0888927
R696 iovdd.n16 iovdd.n14 0.0878254
R697 iovdd.n20 iovdd.n19 0.0878254
R698 iovdd.n496 iovdd.n2 0.0776874
R699 iovdd.n422 iovdd.n400 0.0751466
R700 iovdd.n400 iovdd.n398 0.0751466
R701 iovdd.n397 iovdd.n20 0.0732046
R702 iovdd.n399 iovdd.n14 0.0732046
R703 iovdd.n413 iovdd.n412 0.0727627
R704 iovdd.n412 iovdd.n0 0.0709471
R705 iovdd.n496 iovdd.n495 0.0607875
R706 iovdd.n495 iovdd.n494 0.0607875
R707 iovdd.n494 iovdd.n493 0.0607875
R708 iovdd.n493 iovdd.n492 0.0607875
R709 iovdd.n492 iovdd.n491 0.0607875
R710 iovdd.n491 iovdd.n490 0.0607875
R711 iovdd.n476 iovdd.n32 0.0607875
R712 iovdd.n476 iovdd.n475 0.0607875
R713 iovdd.n475 iovdd.n474 0.0607875
R714 iovdd.n82 iovdd.n72 0.0607875
R715 iovdd.n84 iovdd.n82 0.0607875
R716 iovdd.n86 iovdd.n84 0.0607875
R717 iovdd.n461 iovdd.n460 0.0607875
R718 iovdd.n460 iovdd.n459 0.0607875
R719 iovdd.n459 iovdd.n458 0.0607875
R720 iovdd.n454 iovdd.n453 0.0607875
R721 iovdd.n453 iovdd.n452 0.0607875
R722 iovdd.n452 iovdd.n451 0.0607875
R723 iovdd.n106 iovdd.n97 0.0607875
R724 iovdd.n108 iovdd.n106 0.0607875
R725 iovdd.n110 iovdd.n108 0.0607875
R726 iovdd.n436 iovdd.n435 0.0607875
R727 iovdd.n435 iovdd.n434 0.0607875
R728 iovdd.n434 iovdd.n433 0.0607875
R729 iovdd.n402 iovdd.n117 0.0607875
R730 iovdd.n404 iovdd.n402 0.0607875
R731 iovdd.n406 iovdd.n404 0.0607875
R732 iovdd.n418 iovdd.n417 0.0607875
R733 iovdd.n417 iovdd.n416 0.0607875
R734 iovdd.n183 iovdd.n177 0.0568704
R735 iovdd.n509 iovdd.n2 0.0540779
R736 iovdd.t0 iovdd.n21 0.0491586
R737 iovdd.t0 iovdd.n13 0.048619
R738 iovdd.n490 iovdd.n31 0.045485
R739 iovdd.n501 iovdd.n32 0.045485
R740 iovdd.n458 iovdd.n457 0.045485
R741 iovdd.n455 iovdd.n454 0.045485
R742 iovdd.n111 iovdd.n110 0.045485
R743 iovdd.n438 iovdd.n436 0.045485
R744 iovdd.n407 iovdd.n406 0.045485
R745 iovdd.n420 iovdd.n418 0.045485
R746 iovdd.n416 iovdd.n415 0.045485
R747 iovdd.n473 iovdd.n72 0.0450485
R748 iovdd iovdd.n512 0.0429819
R749 iovdd.n462 iovdd.n86 0.0424295
R750 iovdd.n15 iovdd 0.0411071
R751 iovdd.n451 iovdd.n450 0.0354454
R752 iovdd.n432 iovdd.n117 0.0328263
R753 iovdd.n75 iovdd.t14 0.0323352
R754 iovdd.n19 iovdd.n18 0.0301825
R755 iovdd.n433 iovdd.n432 0.0284612
R756 iovdd.n502 iovdd.n501 0.026254
R757 iovdd.n450 iovdd.n97 0.0258422
R758 iovdd.n18 iovdd 0.0258175
R759 iovdd.n457 iovdd.n91 0.0236349
R760 iovdd.n421 iovdd.n420 0.0210159
R761 iovdd.n462 iovdd.n461 0.0188581
R762 iovdd.n413 iovdd.n394 0.0175238
R763 iovdd.n512 iovdd.n0 0.0169094
R764 iovdd.n439 iovdd.n111 0.0166508
R765 iovdd.n474 iovdd.n473 0.016239
R766 iovdd.n16 iovdd.n15 0.0157896
R767 iovdd.n439 iovdd.n438 0.0140317
R768 iovdd.n415 iovdd.n394 0.0131587
R769 iovdd.n421 iovdd.n407 0.00966667
R770 iovdd.n301 iovdd.n75 0.00930884
R771 iovdd.n190 iovdd.n189 0.00740196
R772 iovdd.n190 iovdd.n172 0.00740196
R773 iovdd.n203 iovdd.n172 0.00740196
R774 iovdd.n204 iovdd.n203 0.00740196
R775 iovdd.n205 iovdd.n204 0.00740196
R776 iovdd.n205 iovdd.n163 0.00740196
R777 iovdd.n218 iovdd.n163 0.00740196
R778 iovdd.n219 iovdd.n218 0.00740196
R779 iovdd.n220 iovdd.n219 0.00740196
R780 iovdd.n220 iovdd.n154 0.00740196
R781 iovdd.n233 iovdd.n154 0.00740196
R782 iovdd.n234 iovdd.n233 0.00740196
R783 iovdd.n260 iovdd.n145 0.00740196
R784 iovdd.n282 iovdd.n281 0.00740196
R785 iovdd.n308 iovdd.n132 0.00740196
R786 iovdd.n390 iovdd.n122 0.00740196
R787 iovdd.n320 iovdd.n122 0.00740196
R788 iovdd.n321 iovdd.n320 0.00740196
R789 iovdd.n329 iovdd.n321 0.00740196
R790 iovdd.n330 iovdd.n329 0.00740196
R791 iovdd.n331 iovdd.n330 0.00740196
R792 iovdd.n339 iovdd.n331 0.00740196
R793 iovdd.n340 iovdd.n339 0.00740196
R794 iovdd.n341 iovdd.n340 0.00740196
R795 iovdd.n349 iovdd.n341 0.00740196
R796 iovdd.n350 iovdd.n349 0.00740196
R797 iovdd.n187 iovdd.n180 0.00740196
R798 iovdd.n191 iovdd.n180 0.00740196
R799 iovdd.n191 iovdd.n173 0.00740196
R800 iovdd.n202 iovdd.n173 0.00740196
R801 iovdd.n202 iovdd.n171 0.00740196
R802 iovdd.n206 iovdd.n171 0.00740196
R803 iovdd.n206 iovdd.n164 0.00740196
R804 iovdd.n217 iovdd.n164 0.00740196
R805 iovdd.n217 iovdd.n162 0.00740196
R806 iovdd.n221 iovdd.n162 0.00740196
R807 iovdd.n221 iovdd.n155 0.00740196
R808 iovdd.n232 iovdd.n155 0.00740196
R809 iovdd.n232 iovdd.n153 0.00740196
R810 iovdd.n248 iovdd.n153 0.00740196
R811 iovdd.n248 iovdd.n146 0.00740196
R812 iovdd.n259 iovdd.n146 0.00740196
R813 iovdd.n259 iovdd.n142 0.00740196
R814 iovdd.n283 iovdd.n142 0.00740196
R815 iovdd.n283 iovdd.n135 0.00740196
R816 iovdd.n294 iovdd.n135 0.00740196
R817 iovdd.n294 iovdd.n131 0.00740196
R818 iovdd.n309 iovdd.n131 0.00740196
R819 iovdd.n309 iovdd.n123 0.00740196
R820 iovdd.n389 iovdd.n123 0.00740196
R821 iovdd.n389 iovdd.n124 0.00740196
R822 iovdd.n382 iovdd.n124 0.00740196
R823 iovdd.n382 iovdd.n381 0.00740196
R824 iovdd.n381 iovdd.n322 0.00740196
R825 iovdd.n374 iovdd.n322 0.00740196
R826 iovdd.n374 iovdd.n373 0.00740196
R827 iovdd.n373 iovdd.n332 0.00740196
R828 iovdd.n366 iovdd.n332 0.00740196
R829 iovdd.n366 iovdd.n365 0.00740196
R830 iovdd.n365 iovdd.n342 0.00740196
R831 iovdd.n358 iovdd.n342 0.00740196
R832 iovdd.n358 iovdd.n357 0.00740196
R833 iovdd.n455 iovdd.n91 0.00704762
R834 iovdd.n247 iovdd.n235 0.00676353
R835 iovdd.n261 iovdd.n143 0.00662549
R836 iovdd.n295 iovdd.n134 0.00648745
R837 iovdd.n307 iovdd.n121 0.00634941
R838 iovdd.n391 iovdd.n121 0.00507255
R839 iovdd.n296 iovdd.n295 0.00493451
R840 iovdd.n280 iovdd.n143 0.00479647
R841 iovdd.n247 iovdd.n246 0.00465843
R842 iovdd.n502 iovdd.n31 0.00442857
R843 iovdd.n357 iovdd.n351 0.00442211
R844 iovdd.n188 iovdd.n187 0.00442211
R845 iovdd.n119 iovdd.n75 0.00437583
R846 iovdd.n186 iovdd.n181 0.00395098
R847 iovdd.n186 iovdd.n185 0.00395098
R848 iovdd.n185 iovdd.n182 0.00395098
R849 iovdd.n182 iovdd.n179 0.00395098
R850 iovdd.n192 iovdd.n179 0.00395098
R851 iovdd.n194 iovdd.n192 0.00395098
R852 iovdd.n194 iovdd.n193 0.00395098
R853 iovdd.n193 iovdd.n174 0.00395098
R854 iovdd.n201 iovdd.n174 0.00395098
R855 iovdd.n201 iovdd.n200 0.00395098
R856 iovdd.n200 iovdd.n175 0.00395098
R857 iovdd.n175 iovdd.n170 0.00395098
R858 iovdd.n207 iovdd.n170 0.00395098
R859 iovdd.n209 iovdd.n207 0.00395098
R860 iovdd.n209 iovdd.n208 0.00395098
R861 iovdd.n208 iovdd.n165 0.00395098
R862 iovdd.n216 iovdd.n165 0.00395098
R863 iovdd.n216 iovdd.n215 0.00395098
R864 iovdd.n215 iovdd.n166 0.00395098
R865 iovdd.n166 iovdd.n161 0.00395098
R866 iovdd.n222 iovdd.n161 0.00395098
R867 iovdd.n224 iovdd.n222 0.00395098
R868 iovdd.n224 iovdd.n223 0.00395098
R869 iovdd.n223 iovdd.n156 0.00395098
R870 iovdd.n231 iovdd.n156 0.00395098
R871 iovdd.n231 iovdd.n230 0.00395098
R872 iovdd.n230 iovdd.n157 0.00395098
R873 iovdd.n157 iovdd.n152 0.00395098
R874 iovdd.n249 iovdd.n152 0.00395098
R875 iovdd.n251 iovdd.n249 0.00395098
R876 iovdd.n251 iovdd.n250 0.00395098
R877 iovdd.n250 iovdd.n147 0.00395098
R878 iovdd.n258 iovdd.n147 0.00395098
R879 iovdd.n258 iovdd.n257 0.00395098
R880 iovdd.n257 iovdd.n148 0.00395098
R881 iovdd.n148 iovdd.n141 0.00395098
R882 iovdd.n284 iovdd.n141 0.00395098
R883 iovdd.n286 iovdd.n284 0.00395098
R884 iovdd.n286 iovdd.n285 0.00395098
R885 iovdd.n285 iovdd.n136 0.00395098
R886 iovdd.n293 iovdd.n136 0.00395098
R887 iovdd.n293 iovdd.n292 0.00395098
R888 iovdd.n292 iovdd.n137 0.00395098
R889 iovdd.n137 iovdd.n130 0.00395098
R890 iovdd.n310 iovdd.n130 0.00395098
R891 iovdd.n312 iovdd.n310 0.00395098
R892 iovdd.n312 iovdd.n311 0.00395098
R893 iovdd.n311 iovdd.n125 0.00395098
R894 iovdd.n388 iovdd.n125 0.00395098
R895 iovdd.n388 iovdd.n387 0.00395098
R896 iovdd.n387 iovdd.n126 0.00395098
R897 iovdd.n384 iovdd.n126 0.00395098
R898 iovdd.n384 iovdd.n383 0.00395098
R899 iovdd.n383 iovdd.n319 0.00395098
R900 iovdd.n380 iovdd.n319 0.00395098
R901 iovdd.n380 iovdd.n379 0.00395098
R902 iovdd.n379 iovdd.n323 0.00395098
R903 iovdd.n376 iovdd.n323 0.00395098
R904 iovdd.n376 iovdd.n375 0.00395098
R905 iovdd.n375 iovdd.n328 0.00395098
R906 iovdd.n372 iovdd.n328 0.00395098
R907 iovdd.n372 iovdd.n371 0.00395098
R908 iovdd.n371 iovdd.n333 0.00395098
R909 iovdd.n368 iovdd.n333 0.00395098
R910 iovdd.n368 iovdd.n367 0.00395098
R911 iovdd.n367 iovdd.n338 0.00395098
R912 iovdd.n364 iovdd.n338 0.00395098
R913 iovdd.n364 iovdd.n363 0.00395098
R914 iovdd.n363 iovdd.n343 0.00395098
R915 iovdd.n360 iovdd.n343 0.00395098
R916 iovdd.n360 iovdd.n359 0.00395098
R917 iovdd.n359 iovdd.n348 0.00395098
R918 iovdd.n356 iovdd.n348 0.00395098
R919 iovdd.n356 iovdd.n355 0.00395098
R920 iovdd.n246 iovdd.n145 0.00324353
R921 iovdd.n282 iovdd.n280 0.00310549
R922 iovdd.n296 iovdd.n132 0.00296745
R923 iovdd.n391 iovdd.n390 0.00282941
R924 iovdd.n354 iovdd 0.00261765
R925 iovdd.n353 iovdd 0.00196667
R926 iovdd.n184 iovdd.n178 0.00191176
R927 iovdd.n195 iovdd.n178 0.00191176
R928 iovdd.n195 iovdd.n176 0.00191176
R929 iovdd.n199 iovdd.n176 0.00191176
R930 iovdd.n199 iovdd.n169 0.00191176
R931 iovdd.n210 iovdd.n169 0.00191176
R932 iovdd.n210 iovdd.n167 0.00191176
R933 iovdd.n214 iovdd.n167 0.00191176
R934 iovdd.n214 iovdd.n160 0.00191176
R935 iovdd.n225 iovdd.n160 0.00191176
R936 iovdd.n225 iovdd.n158 0.00191176
R937 iovdd.n229 iovdd.n158 0.00191176
R938 iovdd.n229 iovdd.n151 0.00191176
R939 iovdd.n252 iovdd.n151 0.00191176
R940 iovdd.n252 iovdd.n149 0.00191176
R941 iovdd.n256 iovdd.n149 0.00191176
R942 iovdd.n256 iovdd.n140 0.00191176
R943 iovdd.n287 iovdd.n140 0.00191176
R944 iovdd.n287 iovdd.n138 0.00191176
R945 iovdd.n291 iovdd.n138 0.00191176
R946 iovdd.n291 iovdd.n129 0.00191176
R947 iovdd.n313 iovdd.n129 0.00191176
R948 iovdd.n313 iovdd.n127 0.00191176
R949 iovdd.n386 iovdd.n127 0.00191176
R950 iovdd.n386 iovdd.n385 0.00191176
R951 iovdd.n385 iovdd.n318 0.00191176
R952 iovdd.n378 iovdd.n318 0.00191176
R953 iovdd.n378 iovdd.n377 0.00191176
R954 iovdd.n377 iovdd.n327 0.00191176
R955 iovdd.n370 iovdd.n327 0.00191176
R956 iovdd.n370 iovdd.n369 0.00191176
R957 iovdd.n369 iovdd.n337 0.00191176
R958 iovdd.n362 iovdd.n337 0.00191176
R959 iovdd.n362 iovdd.n361 0.00191176
R960 iovdd.n361 iovdd.n347 0.00191176
R961 iovdd.n354 iovdd.n347 0.00191176
R962 iovdd.n497 iovdd.n1 0.00170001
R963 iovdd.n184 iovdd.n183 0.0016983
R964 iovdd.n414 iovdd.n35 0.00166668
R965 iovdd.n308 iovdd.n307 0.00155255
R966 iovdd.n196 iovdd.n177 0.00147778
R967 iovdd.n197 iovdd.n196 0.00147778
R968 iovdd.n198 iovdd.n197 0.00147778
R969 iovdd.n198 iovdd.n168 0.00147778
R970 iovdd.n211 iovdd.n168 0.00147778
R971 iovdd.n212 iovdd.n211 0.00147778
R972 iovdd.n213 iovdd.n212 0.00147778
R973 iovdd.n213 iovdd.n159 0.00147778
R974 iovdd.n226 iovdd.n159 0.00147778
R975 iovdd.n227 iovdd.n226 0.00147778
R976 iovdd.n228 iovdd.n227 0.00147778
R977 iovdd.n228 iovdd.n150 0.00147778
R978 iovdd.n253 iovdd.n150 0.00147778
R979 iovdd.n254 iovdd.n253 0.00147778
R980 iovdd.n255 iovdd.n254 0.00147778
R981 iovdd.n255 iovdd.n139 0.00147778
R982 iovdd.n288 iovdd.n139 0.00147778
R983 iovdd.n289 iovdd.n288 0.00147778
R984 iovdd.n290 iovdd.n289 0.00147778
R985 iovdd.n290 iovdd.n128 0.00147778
R986 iovdd.n314 iovdd.n128 0.00147778
R987 iovdd.n315 iovdd.n314 0.00147778
R988 iovdd.n316 iovdd.n315 0.00147778
R989 iovdd.n317 iovdd.n316 0.00147778
R990 iovdd.n324 iovdd.n317 0.00147778
R991 iovdd.n325 iovdd.n324 0.00147778
R992 iovdd.n326 iovdd.n325 0.00147778
R993 iovdd.n334 iovdd.n326 0.00147778
R994 iovdd.n335 iovdd.n334 0.00147778
R995 iovdd.n336 iovdd.n335 0.00147778
R996 iovdd.n344 iovdd.n336 0.00147778
R997 iovdd.n345 iovdd.n344 0.00147778
R998 iovdd.n346 iovdd.n345 0.00147778
R999 iovdd.n352 iovdd.n346 0.00147778
R1000 iovdd.n353 iovdd.n352 0.00147778
R1001 iovdd.n281 iovdd.n134 0.00141451
R1002 iovdd.n411 iovdd.n35 0.00133329
R1003 iovdd.n511 iovdd.n1 0.00129996
R1004 iovdd.n261 iovdd.n260 0.00127647
R1005 iovdd.n235 iovdd.n234 0.00113843
R1006 iovdd.n237 iovdd.n75 0.00100275
R1007 iovdd.n511 iovdd.n13 0.001
R1008 iovdd.n511 iovdd.n21 0.001
R1009 iovdd.n498 iovdd.n484 0.001
R1010 iovdd.n485 iovdd.n483 0.001
R1011 iovdd.n486 iovdd.n482 0.001
R1012 iovdd.n487 iovdd.n481 0.001
R1013 iovdd.n488 iovdd.n480 0.001
R1014 iovdd.n489 iovdd.n479 0.001
R1015 iovdd.n500 iovdd.n33 0.001
R1016 iovdd.n499 iovdd.n34 0.001
R1017 iovdd.n478 iovdd.n477 0.001
R1018 iovdd.n69 iovdd.n68 0.001
R1019 iovdd.n70 iovdd.n67 0.001
R1020 iovdd.n71 iovdd.n66 0.001
R1021 iovdd.n81 iovdd.n65 0.001
R1022 iovdd.n83 iovdd.n64 0.001
R1023 iovdd.n85 iovdd.n63 0.001
R1024 iovdd.n87 iovdd.n62 0.001
R1025 iovdd.n88 iovdd.n61 0.001
R1026 iovdd.n89 iovdd.n60 0.001
R1027 iovdd.n90 iovdd.n59 0.001
R1028 iovdd.n456 iovdd.n58 0.001
R1029 iovdd.n92 iovdd.n57 0.001
R1030 iovdd.n93 iovdd.n56 0.001
R1031 iovdd.n94 iovdd.n55 0.001
R1032 iovdd.n95 iovdd.n54 0.001
R1033 iovdd.n96 iovdd.n53 0.001
R1034 iovdd.n105 iovdd.n52 0.001
R1035 iovdd.n107 iovdd.n51 0.001
R1036 iovdd.n109 iovdd.n50 0.001
R1037 iovdd.n437 iovdd.n49 0.001
R1038 iovdd.n112 iovdd.n48 0.001
R1039 iovdd.n113 iovdd.n47 0.001
R1040 iovdd.n114 iovdd.n46 0.001
R1041 iovdd.n115 iovdd.n45 0.001
R1042 iovdd.n116 iovdd.n44 0.001
R1043 iovdd.n401 iovdd.n43 0.001
R1044 iovdd.n403 iovdd.n42 0.001
R1045 iovdd.n405 iovdd.n41 0.001
R1046 iovdd.n419 iovdd.n40 0.001
R1047 iovdd.n408 iovdd.n39 0.001
R1048 iovdd.n409 iovdd.n38 0.001
R1049 iovdd.n410 iovdd.n37 0.001
R1050 iovdd.n414 iovdd.n36 0.001
R1051 iovdd.n411 iovdd.n13 0.001
R1052 iovdd.n498 iovdd.n497 0.001
R1053 iovdd.n484 iovdd.n483 0.001
R1054 iovdd.n485 iovdd.n482 0.001
R1055 iovdd.n486 iovdd.n481 0.001
R1056 iovdd.n487 iovdd.n480 0.001
R1057 iovdd.n488 iovdd.n479 0.001
R1058 iovdd.n489 iovdd.n33 0.001
R1059 iovdd.n500 iovdd.n499 0.001
R1060 iovdd.n478 iovdd.n34 0.001
R1061 iovdd.n477 iovdd.n68 0.001
R1062 iovdd.n69 iovdd.n67 0.001
R1063 iovdd.n70 iovdd.n66 0.001
R1064 iovdd.n71 iovdd.n65 0.001
R1065 iovdd.n81 iovdd.n64 0.001
R1066 iovdd.n83 iovdd.n63 0.001
R1067 iovdd.n85 iovdd.n62 0.001
R1068 iovdd.n87 iovdd.n61 0.001
R1069 iovdd.n88 iovdd.n60 0.001
R1070 iovdd.n89 iovdd.n59 0.001
R1071 iovdd.n90 iovdd.n58 0.001
R1072 iovdd.n456 iovdd.n57 0.001
R1073 iovdd.n92 iovdd.n56 0.001
R1074 iovdd.n93 iovdd.n55 0.001
R1075 iovdd.n94 iovdd.n54 0.001
R1076 iovdd.n95 iovdd.n53 0.001
R1077 iovdd.n96 iovdd.n52 0.001
R1078 iovdd.n105 iovdd.n51 0.001
R1079 iovdd.n107 iovdd.n50 0.001
R1080 iovdd.n109 iovdd.n49 0.001
R1081 iovdd.n437 iovdd.n48 0.001
R1082 iovdd.n112 iovdd.n47 0.001
R1083 iovdd.n113 iovdd.n46 0.001
R1084 iovdd.n114 iovdd.n45 0.001
R1085 iovdd.n115 iovdd.n44 0.001
R1086 iovdd.n116 iovdd.n43 0.001
R1087 iovdd.n401 iovdd.n42 0.001
R1088 iovdd.n403 iovdd.n41 0.001
R1089 iovdd.n405 iovdd.n40 0.001
R1090 iovdd.n419 iovdd.n39 0.001
R1091 iovdd.n408 iovdd.n38 0.001
R1092 iovdd.n409 iovdd.n37 0.001
R1093 iovdd.n410 iovdd.n36 0.001
R1094 pad.n251 pad 11.7096
R1095 pad pad.t24 9.64317
R1096 pad.n138 pad.n131 4.52159
R1097 pad.n487 pad.n486 4.52158
R1098 pad.n485 pad.n459 4.5005
R1099 pad.n478 pad.n477 4.5005
R1100 pad.n470 pad.n29 4.5005
R1101 pad.n499 pad.n498 4.5005
R1102 pad.n28 pad.n24 4.5005
R1103 pad.n451 pad.n21 4.5005
R1104 pad.n450 pad.n18 4.5005
R1105 pad.n449 pad.n15 4.5005
R1106 pad.n37 pad.n12 4.5005
R1107 pad.n441 pad.n9 4.5005
R1108 pad.n440 pad.n6 4.5005
R1109 pad.n439 pad.n3 4.5005
R1110 pad.n422 pad.n43 4.5005
R1111 pad.n431 pad.n430 4.5005
R1112 pad.n313 pad.n49 4.5005
R1113 pad.n301 pad.n80 4.5005
R1114 pad.n378 pad.n377 4.5005
R1115 pad.n79 pad.n75 4.5005
R1116 pad.n368 pad.n72 4.5005
R1117 pad.n367 pad.n68 4.5005
R1118 pad.n366 pad.n65 4.5005
R1119 pad.n349 pad.n88 4.5005
R1120 pad.n358 pad.n357 4.5005
R1121 pad.n98 pad.n94 4.5005
R1122 pad.n212 pad.n211 4.5005
R1123 pad.n195 pad.n103 4.5005
R1124 pad.n203 pad.n202 4.5005
R1125 pad.n113 pad.n109 4.5005
R1126 pad.n175 pad.n174 4.5005
R1127 pad.n158 pad.n118 4.5005
R1128 pad.n166 pad.n165 4.5005
R1129 pad.n128 pad.n124 4.5005
R1130 pad.n137 pad.n136 4.5005
R1131 pad.n132 pad.n131 4.5005
R1132 pad.n136 pad.n135 4.5005
R1133 pad.n124 pad.n123 4.5005
R1134 pad.n167 pad.n166 4.5005
R1135 pad.n119 pad.n118 4.5005
R1136 pad.n174 pad.n173 4.5005
R1137 pad.n109 pad.n108 4.5005
R1138 pad.n204 pad.n203 4.5005
R1139 pad.n104 pad.n103 4.5005
R1140 pad.n211 pad.n210 4.5005
R1141 pad.n94 pad.n93 4.5005
R1142 pad.n359 pad.n358 4.5005
R1143 pad.n89 pad.n88 4.5005
R1144 pad.n366 pad.n365 4.5005
R1145 pad.n367 pad.n87 4.5005
R1146 pad.n369 pad.n368 4.5005
R1147 pad.n81 pad.n79 4.5005
R1148 pad.n377 pad.n376 4.5005
R1149 pad.n82 pad.n80 4.5005
R1150 pad.n49 pad.n48 4.5005
R1151 pad.n432 pad.n431 4.5005
R1152 pad.n44 pad.n43 4.5005
R1153 pad.n439 pad.n438 4.5005
R1154 pad.n440 pad.n42 4.5005
R1155 pad.n442 pad.n441 4.5005
R1156 pad.n38 pad.n37 4.5005
R1157 pad.n449 pad.n448 4.5005
R1158 pad.n450 pad.n36 4.5005
R1159 pad.n452 pad.n451 4.5005
R1160 pad.n30 pad.n28 4.5005
R1161 pad.n498 pad.n497 4.5005
R1162 pad.n31 pad.n29 4.5005
R1163 pad.n477 pad.n457 4.5005
R1164 pad.n459 pad.n458 4.5005
R1165 pad.n488 pad.n487 4.5005
R1166 pad.n248 pad.n53 4.47552
R1167 pad.n320 pad.n291 4.47552
R1168 pad.n325 pad.n324 4.47552
R1169 pad.n276 pad.n275 4.47552
R1170 pad.n333 pad.n330 4.47552
R1171 pad.n283 pad.n62 4.47552
R1172 pad.n338 pad.n227 4.47552
R1173 pad.n265 pad.n263 4.47552
R1174 pad.n254 pad.n253 3.07063
R1175 pad.n233 pad.n227 3.07063
R1176 pad.n338 pad.n337 3.07063
R1177 pad.n339 pad.n56 3.07063
R1178 pad.n278 pad.n277 3.0005
R1179 pad.n269 pad.n239 3.0005
R1180 pad.n289 pad.n288 3.0005
R1181 pad.n250 pad.n249 3.0005
R1182 pad.n280 pad.n230 3.0005
R1183 pad.n330 pad.n329 3.0005
R1184 pad.n276 pad.n232 3.0005
R1185 pad.n326 pad.n325 3.0005
R1186 pad.n291 pad.n290 3.0005
R1187 pad.n248 pad.n247 3.0005
R1188 pad.n283 pad.n282 3.0005
R1189 pad.n285 pad.n284 3.0005
R1190 pad.n336 pad.n62 3.0005
R1191 pad.n334 pad.n333 3.0005
R1192 pad.n275 pad.n274 3.0005
R1193 pad.n324 pad.n323 3.0005
R1194 pad.n321 pad.n320 3.0005
R1195 pad.n259 pad.n53 3.0005
R1196 pad.n408 pad.n407 3.0005
R1197 pad.n332 pad.n61 3.0005
R1198 pad.n273 pad.n272 3.0005
R1199 pad.n241 pad.n240 3.0005
R1200 pad.n319 pad.n318 3.0005
R1201 pad.n412 pad.n411 3.0005
R1202 pad.n258 pad.n55 3.0005
R1203 pad.n263 pad.n262 3.0005
R1204 pad.n265 pad.n264 3.0005
R1205 pad.n267 pad.n266 3.0005
R1206 pad.n257 pad.t11 2.31826
R1207 pad.n281 pad.t10 2.31826
R1208 pad.n229 pad.t7 2.31826
R1209 pad.n246 pad.t19 2.31826
R1210 pad.n244 pad.t17 2.31826
R1211 pad.n238 pad.t16 2.31826
R1212 pad.n270 pad.t14 2.31826
R1213 pad.n133 pad.n132 2.20699
R1214 pad.n490 pad.n488 2.2005
R1215 pad.n491 pad.n458 2.2005
R1216 pad.n492 pad.n457 2.2005
R1217 pad.n33 pad.n31 2.2005
R1218 pad.n497 pad.n496 2.2005
R1219 pad.n32 pad.n30 2.2005
R1220 pad.n453 pad.n452 2.2005
R1221 pad.n36 pad.n35 2.2005
R1222 pad.n448 pad.n447 2.2005
R1223 pad.n39 pad.n38 2.2005
R1224 pad.n443 pad.n442 2.2005
R1225 pad.n42 pad.n41 2.2005
R1226 pad.n438 pad.n437 2.2005
R1227 pad.n45 pad.n44 2.2005
R1228 pad.n433 pad.n432 2.2005
R1229 pad.n48 pad.n47 2.2005
R1230 pad.n84 pad.n82 2.2005
R1231 pad.n376 pad.n375 2.2005
R1232 pad.n83 pad.n81 2.2005
R1233 pad.n370 pad.n369 2.2005
R1234 pad.n87 pad.n86 2.2005
R1235 pad.n365 pad.n364 2.2005
R1236 pad.n90 pad.n89 2.2005
R1237 pad.n360 pad.n359 2.2005
R1238 pad.n93 pad.n92 2.2005
R1239 pad.n210 pad.n209 2.2005
R1240 pad.n105 pad.n104 2.2005
R1241 pad.n205 pad.n204 2.2005
R1242 pad.n108 pad.n107 2.2005
R1243 pad.n173 pad.n172 2.2005
R1244 pad.n120 pad.n119 2.2005
R1245 pad.n168 pad.n167 2.2005
R1246 pad.n123 pad.n122 2.2005
R1247 pad.n135 pad.n134 2.2005
R1248 pad.n413 pad.t0 1.78531
R1249 pad.n317 pad.t6 1.78531
R1250 pad.n296 pad.t23 1.78531
R1251 pad.n271 pad.t3 1.78531
R1252 pad.n331 pad.t5 1.78531
R1253 pad.n406 pad.t1 1.78531
R1254 pad.n0 pad.t4 1.78531
R1255 pad.n340 pad.t2 1.78502
R1256 pad.n484 pad.n460 1.5005
R1257 pad.n483 pad.n482 1.5005
R1258 pad.n481 pad.n461 1.5005
R1259 pad.n480 pad.n479 1.5005
R1260 pad.n476 pad.n462 1.5005
R1261 pad.n475 pad.n474 1.5005
R1262 pad.n473 pad.n463 1.5005
R1263 pad.n472 pad.n471 1.5005
R1264 pad.n469 pad.n464 1.5005
R1265 pad.n468 pad.n467 1.5005
R1266 pad.n466 pad.n465 1.5005
R1267 pad.n27 pad.n26 1.5005
R1268 pad.n501 pad.n500 1.5005
R1269 pad.n502 pad.n25 1.5005
R1270 pad.n504 pad.n503 1.5005
R1271 pad.n505 pad.n23 1.5005
R1272 pad.n507 pad.n506 1.5005
R1273 pad.n508 pad.n22 1.5005
R1274 pad.n510 pad.n509 1.5005
R1275 pad.n511 pad.n20 1.5005
R1276 pad.n513 pad.n512 1.5005
R1277 pad.n514 pad.n19 1.5005
R1278 pad.n516 pad.n515 1.5005
R1279 pad.n517 pad.n17 1.5005
R1280 pad.n519 pad.n518 1.5005
R1281 pad.n520 pad.n16 1.5005
R1282 pad.n522 pad.n521 1.5005
R1283 pad.n523 pad.n14 1.5005
R1284 pad.n525 pad.n524 1.5005
R1285 pad.n526 pad.n13 1.5005
R1286 pad.n528 pad.n527 1.5005
R1287 pad.n529 pad.n11 1.5005
R1288 pad.n531 pad.n530 1.5005
R1289 pad.n532 pad.n10 1.5005
R1290 pad.n534 pad.n533 1.5005
R1291 pad.n535 pad.n8 1.5005
R1292 pad.n537 pad.n536 1.5005
R1293 pad.n538 pad.n7 1.5005
R1294 pad.n540 pad.n539 1.5005
R1295 pad.n541 pad.n5 1.5005
R1296 pad.n543 pad.n542 1.5005
R1297 pad.n544 pad.n4 1.5005
R1298 pad.n546 pad.n545 1.5005
R1299 pad.n547 pad.n2 1.5005
R1300 pad.n549 pad.n548 1.5005
R1301 pad.n416 pad.n1 1.5005
R1302 pad.n418 pad.n417 1.5005
R1303 pad.n419 pad.n415 1.5005
R1304 pad.n421 pad.n420 1.5005
R1305 pad.n423 pad.n414 1.5005
R1306 pad.n425 pad.n424 1.5005
R1307 pad.n426 pad.n51 1.5005
R1308 pad.n429 pad.n428 1.5005
R1309 pad.n52 pad.n50 1.5005
R1310 pad.n309 pad.n308 1.5005
R1311 pad.n311 pad.n310 1.5005
R1312 pad.n312 pad.n293 1.5005
R1313 pad.n315 pad.n314 1.5005
R1314 pad.n307 pad.n292 1.5005
R1315 pad.n306 pad.n305 1.5005
R1316 pad.n304 pad.n294 1.5005
R1317 pad.n303 pad.n302 1.5005
R1318 pad.n300 pad.n295 1.5005
R1319 pad.n299 pad.n298 1.5005
R1320 pad.n78 pad.n77 1.5005
R1321 pad.n379 pad.n378 1.5005
R1322 pad.n380 pad.n76 1.5005
R1323 pad.n382 pad.n381 1.5005
R1324 pad.n383 pad.n74 1.5005
R1325 pad.n385 pad.n384 1.5005
R1326 pad.n387 pad.n73 1.5005
R1327 pad.n389 pad.n388 1.5005
R1328 pad.n390 pad.n71 1.5005
R1329 pad.n392 pad.n391 1.5005
R1330 pad.n393 pad.n69 1.5005
R1331 pad.n395 pad.n394 1.5005
R1332 pad.n396 pad.n67 1.5005
R1333 pad.n398 pad.n397 1.5005
R1334 pad.n399 pad.n66 1.5005
R1335 pad.n401 pad.n400 1.5005
R1336 pad.n402 pad.n64 1.5005
R1337 pad.n404 pad.n403 1.5005
R1338 pad.n343 pad.n63 1.5005
R1339 pad.n345 pad.n344 1.5005
R1340 pad.n346 pad.n342 1.5005
R1341 pad.n348 pad.n347 1.5005
R1342 pad.n350 pad.n341 1.5005
R1343 pad.n352 pad.n351 1.5005
R1344 pad.n353 pad.n96 1.5005
R1345 pad.n356 pad.n355 1.5005
R1346 pad.n226 pad.n95 1.5005
R1347 pad.n225 pad.n224 1.5005
R1348 pad.n223 pad.n97 1.5005
R1349 pad.n222 pad.n221 1.5005
R1350 pad.n220 pad.n219 1.5005
R1351 pad.n218 pad.n99 1.5005
R1352 pad.n217 pad.n216 1.5005
R1353 pad.n215 pad.n100 1.5005
R1354 pad.n214 pad.n213 1.5005
R1355 pad.n102 pad.n101 1.5005
R1356 pad.n192 pad.n191 1.5005
R1357 pad.n194 pad.n193 1.5005
R1358 pad.n196 pad.n190 1.5005
R1359 pad.n198 pad.n197 1.5005
R1360 pad.n199 pad.n111 1.5005
R1361 pad.n201 pad.n200 1.5005
R1362 pad.n189 pad.n110 1.5005
R1363 pad.n188 pad.n187 1.5005
R1364 pad.n186 pad.n112 1.5005
R1365 pad.n185 pad.n184 1.5005
R1366 pad.n183 pad.n182 1.5005
R1367 pad.n181 pad.n114 1.5005
R1368 pad.n180 pad.n179 1.5005
R1369 pad.n178 pad.n115 1.5005
R1370 pad.n177 pad.n176 1.5005
R1371 pad.n117 pad.n116 1.5005
R1372 pad.n154 pad.n153 1.5005
R1373 pad.n155 pad.n152 1.5005
R1374 pad.n157 pad.n156 1.5005
R1375 pad.n159 pad.n151 1.5005
R1376 pad.n161 pad.n160 1.5005
R1377 pad.n162 pad.n126 1.5005
R1378 pad.n164 pad.n163 1.5005
R1379 pad.n150 pad.n125 1.5005
R1380 pad.n149 pad.n148 1.5005
R1381 pad.n147 pad.n127 1.5005
R1382 pad.n146 pad.n145 1.5005
R1383 pad.n144 pad.n143 1.5005
R1384 pad.n142 pad.n129 1.5005
R1385 pad.n141 pad.n140 1.5005
R1386 pad.n139 pad.n130 1.5005
R1387 pad.n413 pad.n412 1.36955
R1388 pad.n319 pad.n317 1.36955
R1389 pad.n296 pad.n241 1.36955
R1390 pad.n273 pad.n271 1.36955
R1391 pad.n332 pad.n331 1.36955
R1392 pad.n407 pad.n406 1.36955
R1393 pad.n340 pad.n339 1.36955
R1394 pad.n258 pad.n0 1.36955
R1395 pad.n257 pad.t12 1.294
R1396 pad.n281 pad.t13 1.294
R1397 pad.n229 pad.t9 1.294
R1398 pad.n246 pad.t20 1.294
R1399 pad.n244 pad.t8 1.294
R1400 pad.n238 pad.t18 1.294
R1401 pad.n270 pad.t15 1.294
R1402 pad.n251 pad.t21 1.29365
R1403 pad.n252 pad.t22 1.29365
R1404 pad.n122 pad.n121 1.1005
R1405 pad.n169 pad.n168 1.1005
R1406 pad.n170 pad.n120 1.1005
R1407 pad.n172 pad.n171 1.1005
R1408 pad.n107 pad.n106 1.1005
R1409 pad.n206 pad.n205 1.1005
R1410 pad.n207 pad.n105 1.1005
R1411 pad.n209 pad.n208 1.1005
R1412 pad.n92 pad.n91 1.1005
R1413 pad.n361 pad.n360 1.1005
R1414 pad.n362 pad.n90 1.1005
R1415 pad.n364 pad.n363 1.1005
R1416 pad.n86 pad.n85 1.1005
R1417 pad.n371 pad.n370 1.1005
R1418 pad.n372 pad.n83 1.1005
R1419 pad.n375 pad.n374 1.1005
R1420 pad.n373 pad.n84 1.1005
R1421 pad.n47 pad.n46 1.1005
R1422 pad.n434 pad.n433 1.1005
R1423 pad.n435 pad.n45 1.1005
R1424 pad.n437 pad.n436 1.1005
R1425 pad.n41 pad.n40 1.1005
R1426 pad.n444 pad.n443 1.1005
R1427 pad.n445 pad.n39 1.1005
R1428 pad.n447 pad.n446 1.1005
R1429 pad.n35 pad.n34 1.1005
R1430 pad.n454 pad.n453 1.1005
R1431 pad.n455 pad.n32 1.1005
R1432 pad.n496 pad.n495 1.1005
R1433 pad.n494 pad.n33 1.1005
R1434 pad.n493 pad.n492 1.1005
R1435 pad.n491 pad.n456 1.1005
R1436 pad.n490 pad.n489 1.1005
R1437 pad.n249 pad 1.09761
R1438 pad.n289 pad 1.09761
R1439 pad.n239 pad 1.09761
R1440 pad.n277 pad 1.09761
R1441 pad.n230 pad 1.09761
R1442 pad.n284 pad 1.09761
R1443 pad.n253 pad 1.09761
R1444 pad.n266 pad 1.09761
R1445 pad.n252 pad.n251 1.02476
R1446 pad.n427 pad 0.83073
R1447 pad pad.n316 0.83073
R1448 pad.n297 pad 0.83073
R1449 pad.n386 pad 0.83073
R1450 pad pad.n70 0.83073
R1451 pad pad.n405 0.83073
R1452 pad.n354 pad 0.83073
R1453 pad pad.n550 0.83073
R1454 pad.n287 pad.t27 0.672378
R1455 pad.t26 pad.n237 0.672378
R1456 pad.n243 pad.t25 0.672378
R1457 pad.t28 pad.n54 0.672378
R1458 pad.n249 pad.n248 0.64968
R1459 pad.n412 pad.n53 0.64968
R1460 pad.n291 pad.n289 0.64968
R1461 pad.n320 pad.n319 0.64968
R1462 pad.n325 pad.n239 0.64968
R1463 pad.n324 pad.n241 0.64968
R1464 pad.n277 pad.n276 0.64968
R1465 pad.n275 pad.n273 0.64968
R1466 pad.n330 pad.n230 0.64968
R1467 pad.n333 pad.n332 0.64968
R1468 pad.n284 pad.n283 0.64968
R1469 pad.n407 pad.n62 0.64968
R1470 pad.n253 pad.n227 0.64968
R1471 pad.n339 pad.n338 0.64968
R1472 pad.n266 pad.n265 0.64968
R1473 pad.n263 pad.n258 0.64968
R1474 pad.t27 pad.n268 0.589365
R1475 pad.t27 pad.n245 0.589365
R1476 pad.t27 pad.n279 0.589365
R1477 pad.t27 pad.n255 0.589365
R1478 pad.t27 pad.n286 0.589365
R1479 pad.t26 pad.n236 0.589365
R1480 pad.t26 pad.n234 0.589365
R1481 pad.t26 pad.n327 0.589365
R1482 pad.n328 pad.t26 0.589365
R1483 pad.t26 pad.n231 0.589365
R1484 pad.n260 pad.t25 0.589365
R1485 pad.n322 pad.t25 0.589365
R1486 pad.n242 pad.t25 0.589365
R1487 pad.n228 pad.t25 0.589365
R1488 pad.n335 pad.t25 0.589365
R1489 pad.n410 pad.t28 0.589365
R1490 pad.t28 pad.n58 0.589365
R1491 pad.t28 pad.n60 0.589365
R1492 pad.t28 pad.n57 0.589365
R1493 pad.t28 pad.n409 0.589365
R1494 pad.n133 pad.n121 0.557177
R1495 pad pad.n246 0.435451
R1496 pad pad.n244 0.435451
R1497 pad pad.n238 0.435451
R1498 pad pad.n270 0.435451
R1499 pad pad.n229 0.435451
R1500 pad pad.n281 0.435451
R1501 pad pad.n252 0.435451
R1502 pad pad.n257 0.435451
R1503 pad.t27 pad.n256 0.419935
R1504 pad.t26 pad.n235 0.419935
R1505 pad.n261 pad.t25 0.419935
R1506 pad.t28 pad.n59 0.419935
R1507 pad.t27 pad.n254 0.32731
R1508 pad.t26 pad.n233 0.32731
R1509 pad.n337 pad.t25 0.32731
R1510 pad.t28 pad.n56 0.32731
R1511 pad pad.n413 0.317156
R1512 pad.n317 pad 0.317156
R1513 pad pad.n296 0.317156
R1514 pad.n271 pad 0.317156
R1515 pad.n331 pad 0.317156
R1516 pad.n406 pad 0.317156
R1517 pad pad.n340 0.317156
R1518 pad pad.n0 0.317156
R1519 pad.n139 pad.n138 0.278474
R1520 pad.n486 pad.n460 0.278376
R1521 pad.n256 pad 0.188225
R1522 pad.n235 pad 0.188225
R1523 pad.n261 pad 0.188225
R1524 pad.n59 pad 0.188225
R1525 pad.n285 pad.n254 0.183954
R1526 pad.n282 pad.n233 0.183954
R1527 pad.n337 pad.n336 0.183954
R1528 pad.n408 pad.n56 0.183954
R1529 pad.n267 pad.n256 0.160165
R1530 pad.n264 pad.n235 0.160165
R1531 pad.n262 pad.n261 0.160165
R1532 pad.n59 pad.n55 0.160165
R1533 pad.n268 pad.n267 0.146012
R1534 pad.n264 pad.n236 0.146012
R1535 pad.n262 pad.n260 0.146012
R1536 pad.n410 pad.n55 0.146012
R1537 pad.n269 pad.n245 0.140121
R1538 pad.n326 pad.n234 0.140121
R1539 pad.n323 pad.n322 0.140121
R1540 pad.n240 pad.n58 0.140121
R1541 pad.n279 pad.n278 0.136629
R1542 pad.n327 pad.n232 0.136629
R1543 pad.n274 pad.n242 0.136629
R1544 pad.n272 pad.n60 0.136629
R1545 pad.n287 pad.n250 0.135252
R1546 pad.n247 pad.n237 0.135252
R1547 pad.n259 pad.n243 0.135252
R1548 pad.n411 pad.n54 0.135252
R1549 pad.n286 pad.n280 0.13379
R1550 pad.n329 pad.n231 0.13379
R1551 pad.n335 pad.n334 0.13379
R1552 pad.n409 pad.n61 0.13379
R1553 pad.n280 pad.n255 0.133137
R1554 pad.n329 pad.n328 0.133137
R1555 pad.n334 pad.n228 0.133137
R1556 pad.n61 pad.n57 0.133137
R1557 pad.n278 pad.n255 0.130298
R1558 pad.n328 pad.n232 0.130298
R1559 pad.n274 pad.n228 0.130298
R1560 pad.n272 pad.n57 0.130298
R1561 pad.n288 pad.n287 0.129894
R1562 pad.n290 pad.n237 0.129894
R1563 pad.n321 pad.n243 0.129894
R1564 pad.n318 pad.n54 0.129894
R1565 pad.n286 pad.n285 0.129645
R1566 pad.n282 pad.n231 0.129645
R1567 pad.n336 pad.n335 0.129645
R1568 pad.n409 pad.n408 0.129645
R1569 pad.n279 pad.n269 0.126806
R1570 pad.n327 pad.n326 0.126806
R1571 pad.n323 pad.n242 0.126806
R1572 pad.n240 pad.n60 0.126806
R1573 pad.n288 pad.n245 0.123314
R1574 pad.n290 pad.n234 0.123314
R1575 pad.n322 pad.n321 0.123314
R1576 pad.n318 pad.n58 0.123314
R1577 pad.n268 pad.n250 0.117423
R1578 pad.n247 pad.n236 0.117423
R1579 pad.n260 pad.n259 0.117423
R1580 pad.n411 pad.n410 0.117423
R1581 pad.n136 pad.n131 0.0591667
R1582 pad.n136 pad.n124 0.0591667
R1583 pad.n166 pad.n124 0.0591667
R1584 pad.n166 pad.n118 0.0591667
R1585 pad.n174 pad.n118 0.0591667
R1586 pad.n174 pad.n109 0.0591667
R1587 pad.n203 pad.n109 0.0591667
R1588 pad.n203 pad.n103 0.0591667
R1589 pad.n211 pad.n103 0.0591667
R1590 pad.n211 pad.n94 0.0591667
R1591 pad.n358 pad.n94 0.0591667
R1592 pad.n358 pad.n88 0.0591667
R1593 pad.n366 pad.n88 0.0591667
R1594 pad.n367 pad.n366 0.0591667
R1595 pad.n368 pad.n367 0.0591667
R1596 pad.n368 pad.n79 0.0591667
R1597 pad.n377 pad.n79 0.0591667
R1598 pad.n377 pad.n80 0.0591667
R1599 pad.n80 pad.n49 0.0591667
R1600 pad.n431 pad.n49 0.0591667
R1601 pad.n431 pad.n43 0.0591667
R1602 pad.n439 pad.n43 0.0591667
R1603 pad.n440 pad.n439 0.0591667
R1604 pad.n441 pad.n440 0.0591667
R1605 pad.n441 pad.n37 0.0591667
R1606 pad.n449 pad.n37 0.0591667
R1607 pad.n450 pad.n449 0.0591667
R1608 pad.n451 pad.n450 0.0591667
R1609 pad.n451 pad.n28 0.0591667
R1610 pad.n498 pad.n28 0.0591667
R1611 pad.n498 pad.n29 0.0591667
R1612 pad.n477 pad.n29 0.0591667
R1613 pad.n477 pad.n459 0.0591667
R1614 pad.n487 pad.n459 0.0591667
R1615 pad.n135 pad.n132 0.0591667
R1616 pad.n135 pad.n123 0.0591667
R1617 pad.n167 pad.n123 0.0591667
R1618 pad.n167 pad.n119 0.0591667
R1619 pad.n173 pad.n119 0.0591667
R1620 pad.n173 pad.n108 0.0591667
R1621 pad.n204 pad.n108 0.0591667
R1622 pad.n204 pad.n104 0.0591667
R1623 pad.n210 pad.n104 0.0591667
R1624 pad.n210 pad.n93 0.0591667
R1625 pad.n359 pad.n93 0.0591667
R1626 pad.n359 pad.n89 0.0591667
R1627 pad.n365 pad.n89 0.0591667
R1628 pad.n365 pad.n87 0.0591667
R1629 pad.n369 pad.n87 0.0591667
R1630 pad.n369 pad.n81 0.0591667
R1631 pad.n376 pad.n81 0.0591667
R1632 pad.n376 pad.n82 0.0591667
R1633 pad.n82 pad.n48 0.0591667
R1634 pad.n432 pad.n48 0.0591667
R1635 pad.n432 pad.n44 0.0591667
R1636 pad.n438 pad.n44 0.0591667
R1637 pad.n438 pad.n42 0.0591667
R1638 pad.n442 pad.n42 0.0591667
R1639 pad.n442 pad.n38 0.0591667
R1640 pad.n448 pad.n38 0.0591667
R1641 pad.n448 pad.n36 0.0591667
R1642 pad.n452 pad.n36 0.0591667
R1643 pad.n452 pad.n30 0.0591667
R1644 pad.n497 pad.n30 0.0591667
R1645 pad.n497 pad.n31 0.0591667
R1646 pad.n457 pad.n31 0.0591667
R1647 pad.n458 pad.n457 0.0591667
R1648 pad.n488 pad.n458 0.0591667
R1649 pad.n486 pad.n485 0.0407494
R1650 pad.n138 pad.n137 0.0407425
R1651 pad.n140 pad.n139 0.0148733
R1652 pad.n140 pad.n129 0.0148733
R1653 pad.n144 pad.n129 0.0148733
R1654 pad.n145 pad.n144 0.0148733
R1655 pad.n145 pad.n127 0.0148733
R1656 pad.n149 pad.n127 0.0148733
R1657 pad.n150 pad.n149 0.0148733
R1658 pad.n163 pad.n150 0.0148733
R1659 pad.n163 pad.n162 0.0148733
R1660 pad.n162 pad.n161 0.0148733
R1661 pad.n161 pad.n151 0.0148733
R1662 pad.n156 pad.n151 0.0148733
R1663 pad.n156 pad.n155 0.0148733
R1664 pad.n155 pad.n154 0.0148733
R1665 pad.n154 pad.n116 0.0148733
R1666 pad.n177 pad.n116 0.0148733
R1667 pad.n178 pad.n177 0.0148733
R1668 pad.n179 pad.n178 0.0148733
R1669 pad.n179 pad.n114 0.0148733
R1670 pad.n183 pad.n114 0.0148733
R1671 pad.n184 pad.n183 0.0148733
R1672 pad.n184 pad.n112 0.0148733
R1673 pad.n188 pad.n112 0.0148733
R1674 pad.n189 pad.n188 0.0148733
R1675 pad.n200 pad.n189 0.0148733
R1676 pad.n200 pad.n199 0.0148733
R1677 pad.n199 pad.n198 0.0148733
R1678 pad.n198 pad.n190 0.0148733
R1679 pad.n193 pad.n190 0.0148733
R1680 pad.n193 pad.n192 0.0148733
R1681 pad.n192 pad.n101 0.0148733
R1682 pad.n214 pad.n101 0.0148733
R1683 pad.n215 pad.n214 0.0148733
R1684 pad.n216 pad.n215 0.0148733
R1685 pad.n216 pad.n99 0.0148733
R1686 pad.n220 pad.n99 0.0148733
R1687 pad.n221 pad.n220 0.0148733
R1688 pad.n221 pad.n97 0.0148733
R1689 pad.n225 pad.n97 0.0148733
R1690 pad.n226 pad.n225 0.0148733
R1691 pad.n355 pad.n226 0.0148733
R1692 pad.n353 pad.n352 0.0148733
R1693 pad.n352 pad.n341 0.0148733
R1694 pad.n347 pad.n341 0.0148733
R1695 pad.n347 pad.n346 0.0148733
R1696 pad.n346 pad.n345 0.0148733
R1697 pad.n345 pad.n63 0.0148733
R1698 pad.n404 pad.n64 0.0148733
R1699 pad.n400 pad.n64 0.0148733
R1700 pad.n400 pad.n399 0.0148733
R1701 pad.n399 pad.n398 0.0148733
R1702 pad.n398 pad.n67 0.0148733
R1703 pad.n394 pad.n393 0.0148733
R1704 pad.n393 pad.n392 0.0148733
R1705 pad.n392 pad.n71 0.0148733
R1706 pad.n388 pad.n71 0.0148733
R1707 pad.n388 pad.n387 0.0148733
R1708 pad.n385 pad.n74 0.0148733
R1709 pad.n381 pad.n74 0.0148733
R1710 pad.n381 pad.n380 0.0148733
R1711 pad.n380 pad.n379 0.0148733
R1712 pad.n379 pad.n77 0.0148733
R1713 pad.n298 pad.n295 0.0148733
R1714 pad.n303 pad.n295 0.0148733
R1715 pad.n304 pad.n303 0.0148733
R1716 pad.n305 pad.n304 0.0148733
R1717 pad.n305 pad.n292 0.0148733
R1718 pad.n315 pad.n293 0.0148733
R1719 pad.n310 pad.n293 0.0148733
R1720 pad.n310 pad.n309 0.0148733
R1721 pad.n309 pad.n52 0.0148733
R1722 pad.n428 pad.n52 0.0148733
R1723 pad.n426 pad.n425 0.0148733
R1724 pad.n425 pad.n414 0.0148733
R1725 pad.n420 pad.n414 0.0148733
R1726 pad.n420 pad.n419 0.0148733
R1727 pad.n419 pad.n418 0.0148733
R1728 pad.n418 pad.n1 0.0148733
R1729 pad.n549 pad.n2 0.0148733
R1730 pad.n545 pad.n2 0.0148733
R1731 pad.n545 pad.n544 0.0148733
R1732 pad.n544 pad.n543 0.0148733
R1733 pad.n543 pad.n5 0.0148733
R1734 pad.n539 pad.n5 0.0148733
R1735 pad.n539 pad.n538 0.0148733
R1736 pad.n538 pad.n537 0.0148733
R1737 pad.n537 pad.n8 0.0148733
R1738 pad.n533 pad.n8 0.0148733
R1739 pad.n533 pad.n532 0.0148733
R1740 pad.n532 pad.n531 0.0148733
R1741 pad.n531 pad.n11 0.0148733
R1742 pad.n527 pad.n11 0.0148733
R1743 pad.n527 pad.n526 0.0148733
R1744 pad.n526 pad.n525 0.0148733
R1745 pad.n525 pad.n14 0.0148733
R1746 pad.n521 pad.n14 0.0148733
R1747 pad.n521 pad.n520 0.0148733
R1748 pad.n520 pad.n519 0.0148733
R1749 pad.n519 pad.n17 0.0148733
R1750 pad.n515 pad.n17 0.0148733
R1751 pad.n515 pad.n514 0.0148733
R1752 pad.n514 pad.n513 0.0148733
R1753 pad.n513 pad.n20 0.0148733
R1754 pad.n509 pad.n20 0.0148733
R1755 pad.n509 pad.n508 0.0148733
R1756 pad.n508 pad.n507 0.0148733
R1757 pad.n507 pad.n23 0.0148733
R1758 pad.n503 pad.n23 0.0148733
R1759 pad.n503 pad.n502 0.0148733
R1760 pad.n502 pad.n501 0.0148733
R1761 pad.n501 pad.n26 0.0148733
R1762 pad.n466 pad.n26 0.0148733
R1763 pad.n467 pad.n466 0.0148733
R1764 pad.n467 pad.n464 0.0148733
R1765 pad.n472 pad.n464 0.0148733
R1766 pad.n473 pad.n472 0.0148733
R1767 pad.n474 pad.n473 0.0148733
R1768 pad.n474 pad.n462 0.0148733
R1769 pad.n480 pad.n462 0.0148733
R1770 pad.n481 pad.n480 0.0148733
R1771 pad.n482 pad.n481 0.0148733
R1772 pad.n482 pad.n460 0.0148733
R1773 pad.n141 pad.n130 0.0148733
R1774 pad.n142 pad.n141 0.0148733
R1775 pad.n143 pad.n142 0.0148733
R1776 pad.n147 pad.n146 0.0148733
R1777 pad.n148 pad.n147 0.0148733
R1778 pad.n148 pad.n125 0.0148733
R1779 pad.n164 pad.n126 0.0148733
R1780 pad.n160 pad.n126 0.0148733
R1781 pad.n160 pad.n159 0.0148733
R1782 pad.n157 pad.n152 0.0148733
R1783 pad.n153 pad.n152 0.0148733
R1784 pad.n153 pad.n117 0.0148733
R1785 pad.n176 pad.n117 0.0148733
R1786 pad.n180 pad.n115 0.0148733
R1787 pad.n181 pad.n180 0.0148733
R1788 pad.n182 pad.n181 0.0148733
R1789 pad.n186 pad.n185 0.0148733
R1790 pad.n187 pad.n186 0.0148733
R1791 pad.n187 pad.n110 0.0148733
R1792 pad.n201 pad.n111 0.0148733
R1793 pad.n197 pad.n111 0.0148733
R1794 pad.n197 pad.n196 0.0148733
R1795 pad.n194 pad.n191 0.0148733
R1796 pad.n191 pad.n102 0.0148733
R1797 pad.n213 pad.n102 0.0148733
R1798 pad.n217 pad.n100 0.0148733
R1799 pad.n218 pad.n217 0.0148733
R1800 pad.n219 pad.n218 0.0148733
R1801 pad.n223 pad.n222 0.0148733
R1802 pad.n224 pad.n223 0.0148733
R1803 pad.n224 pad.n95 0.0148733
R1804 pad.n356 pad.n96 0.0148733
R1805 pad.n351 pad.n96 0.0148733
R1806 pad.n351 pad.n350 0.0148733
R1807 pad.n348 pad.n342 0.0148733
R1808 pad.n344 pad.n342 0.0148733
R1809 pad.n344 pad.n343 0.0148733
R1810 pad.n403 pad.n402 0.0148733
R1811 pad.n402 pad.n401 0.0148733
R1812 pad.n401 pad.n66 0.0148733
R1813 pad.n397 pad.n396 0.0148733
R1814 pad.n396 pad.n395 0.0148733
R1815 pad.n395 pad.n69 0.0148733
R1816 pad.n391 pad.n390 0.0148733
R1817 pad.n390 pad.n389 0.0148733
R1818 pad.n389 pad.n73 0.0148733
R1819 pad.n384 pad.n383 0.0148733
R1820 pad.n383 pad.n382 0.0148733
R1821 pad.n382 pad.n76 0.0148733
R1822 pad.n378 pad.n76 0.0148733
R1823 pad.n378 pad.n78 0.0148733
R1824 pad.n299 pad.n78 0.0148733
R1825 pad.n300 pad.n299 0.0148733
R1826 pad.n302 pad.n300 0.0148733
R1827 pad.n306 pad.n294 0.0148733
R1828 pad.n307 pad.n306 0.0148733
R1829 pad.n314 pad.n307 0.0148733
R1830 pad.n312 pad.n311 0.0148733
R1831 pad.n311 pad.n308 0.0148733
R1832 pad.n308 pad.n50 0.0148733
R1833 pad.n429 pad.n51 0.0148733
R1834 pad.n424 pad.n51 0.0148733
R1835 pad.n424 pad.n423 0.0148733
R1836 pad.n421 pad.n415 0.0148733
R1837 pad.n417 pad.n415 0.0148733
R1838 pad.n417 pad.n416 0.0148733
R1839 pad.n548 pad.n547 0.0148733
R1840 pad.n547 pad.n546 0.0148733
R1841 pad.n546 pad.n4 0.0148733
R1842 pad.n542 pad.n541 0.0148733
R1843 pad.n541 pad.n540 0.0148733
R1844 pad.n540 pad.n7 0.0148733
R1845 pad.n536 pad.n535 0.0148733
R1846 pad.n535 pad.n534 0.0148733
R1847 pad.n534 pad.n10 0.0148733
R1848 pad.n530 pad.n529 0.0148733
R1849 pad.n529 pad.n528 0.0148733
R1850 pad.n528 pad.n13 0.0148733
R1851 pad.n524 pad.n523 0.0148733
R1852 pad.n523 pad.n522 0.0148733
R1853 pad.n522 pad.n16 0.0148733
R1854 pad.n518 pad.n517 0.0148733
R1855 pad.n517 pad.n516 0.0148733
R1856 pad.n516 pad.n19 0.0148733
R1857 pad.n512 pad.n511 0.0148733
R1858 pad.n511 pad.n510 0.0148733
R1859 pad.n510 pad.n22 0.0148733
R1860 pad.n506 pad.n505 0.0148733
R1861 pad.n505 pad.n504 0.0148733
R1862 pad.n504 pad.n25 0.0148733
R1863 pad.n500 pad.n25 0.0148733
R1864 pad.n465 pad.n27 0.0148733
R1865 pad.n468 pad.n465 0.0148733
R1866 pad.n469 pad.n468 0.0148733
R1867 pad.n471 pad.n463 0.0148733
R1868 pad.n475 pad.n463 0.0148733
R1869 pad.n476 pad.n475 0.0148733
R1870 pad.n479 pad.n461 0.0148733
R1871 pad.n483 pad.n461 0.0148733
R1872 pad.n484 pad.n483 0.0148733
R1873 pad.n175 pad.n115 0.01458
R1874 pad.n24 pad.n22 0.01458
R1875 pad.n550 pad.n549 0.0144333
R1876 pad.n405 pad.n404 0.01414
R1877 pad.n159 pad.n158 0.0139933
R1878 pad.n499 pad.n27 0.0139933
R1879 pad.n75 pad.n73 0.0137
R1880 pad.n301 pad.n294 0.0137
R1881 pad.n185 pad.n113 0.0134067
R1882 pad.n21 pad.n19 0.0134067
R1883 pad.n355 pad.n354 0.01326
R1884 pad.n428 pad.n427 0.0129667
R1885 pad.n165 pad.n125 0.01282
R1886 pad.n471 pad.n470 0.01282
R1887 pad.n72 pad.n69 0.0125267
R1888 pad.n313 pad.n312 0.0125267
R1889 pad.n134 pad.n122 0.0125
R1890 pad.n168 pad.n122 0.0125
R1891 pad.n168 pad.n120 0.0125
R1892 pad.n172 pad.n120 0.0125
R1893 pad.n172 pad.n107 0.0125
R1894 pad.n205 pad.n107 0.0125
R1895 pad.n205 pad.n105 0.0125
R1896 pad.n209 pad.n105 0.0125
R1897 pad.n209 pad.n92 0.0125
R1898 pad.n360 pad.n92 0.0125
R1899 pad.n360 pad.n90 0.0125
R1900 pad.n364 pad.n90 0.0125
R1901 pad.n364 pad.n86 0.0125
R1902 pad.n370 pad.n86 0.0125
R1903 pad.n370 pad.n83 0.0125
R1904 pad.n375 pad.n83 0.0125
R1905 pad.n375 pad.n84 0.0125
R1906 pad.n84 pad.n47 0.0125
R1907 pad.n433 pad.n47 0.0125
R1908 pad.n433 pad.n45 0.0125
R1909 pad.n437 pad.n45 0.0125
R1910 pad.n437 pad.n41 0.0125
R1911 pad.n443 pad.n41 0.0125
R1912 pad.n443 pad.n39 0.0125
R1913 pad.n447 pad.n39 0.0125
R1914 pad.n447 pad.n35 0.0125
R1915 pad.n453 pad.n35 0.0125
R1916 pad.n453 pad.n32 0.0125
R1917 pad.n496 pad.n32 0.0125
R1918 pad.n496 pad.n33 0.0125
R1919 pad.n492 pad.n33 0.0125
R1920 pad.n492 pad.n491 0.0125
R1921 pad.n491 pad.n490 0.0125
R1922 pad.n202 pad.n201 0.0122333
R1923 pad.n18 pad.n16 0.0122333
R1924 pad.n394 pad.n70 0.0117933
R1925 pad.n143 pad.n128 0.0116467
R1926 pad.n479 pad.n478 0.0116467
R1927 pad.n68 pad.n66 0.0113533
R1928 pad.n430 pad.n429 0.0113533
R1929 pad.n195 pad.n194 0.01106
R1930 pad.n15 pad.n13 0.01106
R1931 pad.n316 pad.n292 0.01062
R1932 pad.n343 pad.n65 0.01018
R1933 pad.n422 pad.n421 0.01018
R1934 pad.n212 pad.n100 0.00988667
R1935 pad.n12 pad.n10 0.00988667
R1936 pad.n386 pad.n385 0.00944667
R1937 pad.n350 pad.n349 0.00900667
R1938 pad.n548 pad.n3 0.00900667
R1939 pad.n222 pad.n98 0.00871333
R1940 pad.n9 pad.n7 0.00871333
R1941 pad.n297 pad.n77 0.00827333
R1942 pad.n357 pad.n95 0.00783333
R1943 pad.n542 pad.n6 0.00783333
R1944 pad.n169 pad.n121 0.00783333
R1945 pad.n170 pad.n169 0.00783333
R1946 pad.n171 pad.n170 0.00783333
R1947 pad.n171 pad.n106 0.00783333
R1948 pad.n206 pad.n106 0.00783333
R1949 pad.n207 pad.n206 0.00783333
R1950 pad.n208 pad.n207 0.00783333
R1951 pad.n208 pad.n91 0.00783333
R1952 pad.n361 pad.n91 0.00783333
R1953 pad.n362 pad.n361 0.00783333
R1954 pad.n363 pad.n362 0.00783333
R1955 pad.n363 pad.n85 0.00783333
R1956 pad.n371 pad.n85 0.00783333
R1957 pad.n372 pad.n371 0.00783333
R1958 pad.n374 pad.n372 0.00783333
R1959 pad.n374 pad.n373 0.00783333
R1960 pad.n373 pad.n46 0.00783333
R1961 pad.n434 pad.n46 0.00783333
R1962 pad.n435 pad.n434 0.00783333
R1963 pad.n436 pad.n435 0.00783333
R1964 pad.n436 pad.n40 0.00783333
R1965 pad.n444 pad.n40 0.00783333
R1966 pad.n445 pad.n444 0.00783333
R1967 pad.n446 pad.n445 0.00783333
R1968 pad.n446 pad.n34 0.00783333
R1969 pad.n454 pad.n34 0.00783333
R1970 pad.n455 pad.n454 0.00783333
R1971 pad.n495 pad.n455 0.00783333
R1972 pad.n495 pad.n494 0.00783333
R1973 pad.n494 pad.n493 0.00783333
R1974 pad.n493 pad.n456 0.00783333
R1975 pad.n489 pad.n456 0.00783333
R1976 pad.n357 pad.n356 0.00754
R1977 pad.n6 pad.n4 0.00754
R1978 pad.n298 pad.n297 0.0071
R1979 pad.n134 pad.n133 0.00694773
R1980 pad.n219 pad.n98 0.00666
R1981 pad.n536 pad.n9 0.00666
R1982 pad.n349 pad.n348 0.00636667
R1983 pad.n416 pad.n3 0.00636667
R1984 pad.n387 pad.n386 0.00592667
R1985 pad.n213 pad.n212 0.00548667
R1986 pad.n530 pad.n12 0.00548667
R1987 pad.n403 pad.n65 0.00519333
R1988 pad.n423 pad.n422 0.00519333
R1989 pad.n137 pad.n130 0.0049
R1990 pad.n485 pad.n484 0.0049
R1991 pad.n316 pad.n315 0.00475333
R1992 pad.n196 pad.n195 0.00431333
R1993 pad.n524 pad.n15 0.00431333
R1994 pad.n489 pad 0.00416667
R1995 pad.n397 pad.n68 0.00402
R1996 pad.n430 pad.n50 0.00402
R1997 pad.n146 pad.n128 0.00372667
R1998 pad.n478 pad.n476 0.00372667
R1999 pad.n70 pad.n67 0.00358
R2000 pad.n202 pad.n110 0.00314
R2001 pad.n518 pad.n18 0.00314
R2002 pad.n391 pad.n72 0.00284667
R2003 pad.n314 pad.n313 0.00284667
R2004 pad.n165 pad.n164 0.00255333
R2005 pad.n470 pad.n469 0.00255333
R2006 pad.n427 pad.n426 0.00240667
R2007 pad.n354 pad.n353 0.00211333
R2008 pad.n182 pad.n113 0.00196667
R2009 pad.n512 pad.n21 0.00196667
R2010 pad.n384 pad.n75 0.00167333
R2011 pad.n302 pad.n301 0.00167333
R2012 pad.n158 pad.n157 0.00138
R2013 pad.n500 pad.n499 0.00138
R2014 pad.n405 pad.n63 0.00123333
R2015 pad.n550 pad.n1 0.00094
R2016 pad.n176 pad.n175 0.000793333
R2017 pad.n506 pad.n24 0.000793333
R2018 sg13g2_GateDecode_0.sg13g2_LevelUp_0.o sg13g2_Clamp_N15N15D_0.gate 60.0387
R2019 sg13g2_GateDecode_0.ngate.n15 sg13g2_GateDecode_0.ngate.n14 9.75711
R2020 sg13g2_GateDecode_0.ngate.n1 sg13g2_GateDecode_0.ngate.t3 9.10182
R2021 sg13g2_GateDecode_0.ngate.n13 sg13g2_GateDecode_0.ngate.t2 8.24932
R2022 sg13g2_GateDecode_0.ngate.n12 sg13g2_GateDecode_0.ngate.t7 8.24932
R2023 sg13g2_GateDecode_0.ngate.n11 sg13g2_GateDecode_0.ngate.t13 8.24932
R2024 sg13g2_GateDecode_0.ngate.n10 sg13g2_GateDecode_0.ngate.t4 8.24932
R2025 sg13g2_GateDecode_0.ngate.n9 sg13g2_GateDecode_0.ngate.t14 8.24932
R2026 sg13g2_GateDecode_0.ngate.n8 sg13g2_GateDecode_0.ngate.t17 8.24932
R2027 sg13g2_GateDecode_0.ngate.n7 sg13g2_GateDecode_0.ngate.t6 8.24932
R2028 sg13g2_GateDecode_0.ngate.n6 sg13g2_GateDecode_0.ngate.t16 8.24932
R2029 sg13g2_GateDecode_0.ngate.n5 sg13g2_GateDecode_0.ngate.t8 8.24932
R2030 sg13g2_GateDecode_0.ngate.n4 sg13g2_GateDecode_0.ngate.t9 8.24932
R2031 sg13g2_GateDecode_0.ngate.n3 sg13g2_GateDecode_0.ngate.t5 8.24932
R2032 sg13g2_GateDecode_0.ngate.n2 sg13g2_GateDecode_0.ngate.t11 8.24932
R2033 sg13g2_GateDecode_0.ngate.n1 sg13g2_GateDecode_0.ngate.t15 8.24932
R2034 sg13g2_GateDecode_0.ngate.n14 sg13g2_GateDecode_0.ngate.t10 8.24932
R2035 sg13g2_GateDecode_0.ngate.n0 sg13g2_GateDecode_0.ngate.t0 4.59834
R2036 sg13g2_GateDecode_0.ngate.n16 sg13g2_GateDecode_0.ngate.n15 4.5005
R2037 sg13g2_GateDecode_0.ngate.n15 sg13g2_GateDecode_0.ngate.t12 4.31293
R2038 sg13g2_GateDecode_0.ngate.n0 sg13g2_GateDecode_0.ngate.t1 2.00385
R2039 sg13g2_GateDecode_0.sg13g2_LevelUp_0.o sg13g2_GateDecode_0.ngate.n0 1.98894
R2040 sg13g2_GateDecode_0.ngate.n2 sg13g2_GateDecode_0.ngate.n1 1.22425
R2041 sg13g2_GateDecode_0.ngate.n4 sg13g2_GateDecode_0.ngate.n3 1.22425
R2042 sg13g2_GateDecode_0.ngate.n6 sg13g2_GateDecode_0.ngate.n5 1.22425
R2043 sg13g2_GateDecode_0.ngate.n8 sg13g2_GateDecode_0.ngate.n7 1.22425
R2044 sg13g2_GateDecode_0.ngate.n10 sg13g2_GateDecode_0.ngate.n9 1.22425
R2045 sg13g2_GateDecode_0.ngate.n12 sg13g2_GateDecode_0.ngate.n11 1.22425
R2046 sg13g2_GateDecode_0.ngate.n14 sg13g2_GateDecode_0.ngate.n13 1.22425
R2047 sg13g2_Clamp_N15N15D_0.gate sg13g2_GateDecode_0.ngate.n16 1.17264
R2048 sg13g2_GateDecode_0.ngate.n3 sg13g2_GateDecode_0.ngate.n2 0.853
R2049 sg13g2_GateDecode_0.ngate.n5 sg13g2_GateDecode_0.ngate.n4 0.853
R2050 sg13g2_GateDecode_0.ngate.n7 sg13g2_GateDecode_0.ngate.n6 0.853
R2051 sg13g2_GateDecode_0.ngate.n9 sg13g2_GateDecode_0.ngate.n8 0.853
R2052 sg13g2_GateDecode_0.ngate.n11 sg13g2_GateDecode_0.ngate.n10 0.853
R2053 sg13g2_GateDecode_0.ngate.n13 sg13g2_GateDecode_0.ngate.n12 0.853
R2054 sg13g2_GateDecode_0.ngate.n16 sg13g2_Clamp_N15N15D_0.gate 0.1545
R2055 iovss.n220 iovss.n219 0.826084
R2056 iovss.n84 iovss.n80 0.826084
R2057 iovss.n218 iovss.n217 0.818682
R2058 iovss.n5 iovss.n4 0.818682
R2059 iovss.n206 iovss.n205 0.818682
R2060 iovss.n204 iovss.n12 0.818682
R2061 iovss.n203 iovss.n202 0.818682
R2062 iovss.n14 iovss.n13 0.818682
R2063 iovss.n191 iovss.n190 0.818682
R2064 iovss.n189 iovss.n21 0.818682
R2065 iovss.n188 iovss.n187 0.818682
R2066 iovss.n23 iovss.n22 0.818682
R2067 iovss.n176 iovss.n175 0.818682
R2068 iovss.n174 iovss.n30 0.818682
R2069 iovss.n173 iovss.n172 0.818682
R2070 iovss.n32 iovss.n31 0.818682
R2071 iovss.n161 iovss.n160 0.818682
R2072 iovss.n159 iovss.n39 0.818682
R2073 iovss.n158 iovss.n157 0.818682
R2074 iovss.n41 iovss.n40 0.818682
R2075 iovss.n146 iovss.n145 0.818682
R2076 iovss.n144 iovss.n48 0.818682
R2077 iovss.n143 iovss.n142 0.818682
R2078 iovss.n50 iovss.n49 0.818682
R2079 iovss.n131 iovss.n130 0.818682
R2080 iovss.n129 iovss.n57 0.818682
R2081 iovss.n128 iovss.n127 0.818682
R2082 iovss.n59 iovss.n58 0.818682
R2083 iovss.n116 iovss.n115 0.818682
R2084 iovss.n114 iovss.n66 0.818682
R2085 iovss.n113 iovss.n112 0.818682
R2086 iovss.n68 iovss.n67 0.818682
R2087 iovss.n101 iovss.n100 0.818682
R2088 iovss.n99 iovss.n75 0.818682
R2089 iovss.n98 iovss.n97 0.818682
R2090 iovss.n77 iovss.n76 0.818682
R2091 iovss.n86 iovss.n85 0.818682
R2092 iovss.n83 iovss.n81 0.818682
R2093 iovss.n87 iovss.n86 0.818682
R2094 iovss.n78 iovss.n77 0.818682
R2095 iovss.n97 iovss.n96 0.818682
R2096 iovss.n75 iovss.n73 0.818682
R2097 iovss.n102 iovss.n101 0.818682
R2098 iovss.n69 iovss.n68 0.818682
R2099 iovss.n112 iovss.n111 0.818682
R2100 iovss.n66 iovss.n64 0.818682
R2101 iovss.n117 iovss.n116 0.818682
R2102 iovss.n60 iovss.n59 0.818682
R2103 iovss.n127 iovss.n126 0.818682
R2104 iovss.n57 iovss.n55 0.818682
R2105 iovss.n132 iovss.n131 0.818682
R2106 iovss.n51 iovss.n50 0.818682
R2107 iovss.n142 iovss.n141 0.818682
R2108 iovss.n48 iovss.n46 0.818682
R2109 iovss.n147 iovss.n146 0.818682
R2110 iovss.n42 iovss.n41 0.818682
R2111 iovss.n157 iovss.n156 0.818682
R2112 iovss.n39 iovss.n37 0.818682
R2113 iovss.n162 iovss.n161 0.818682
R2114 iovss.n33 iovss.n32 0.818682
R2115 iovss.n172 iovss.n171 0.818682
R2116 iovss.n30 iovss.n28 0.818682
R2117 iovss.n177 iovss.n176 0.818682
R2118 iovss.n24 iovss.n23 0.818682
R2119 iovss.n187 iovss.n186 0.818682
R2120 iovss.n21 iovss.n19 0.818682
R2121 iovss.n192 iovss.n191 0.818682
R2122 iovss.n15 iovss.n14 0.818682
R2123 iovss.n202 iovss.n201 0.818682
R2124 iovss.n12 iovss.n10 0.818682
R2125 iovss.n207 iovss.n206 0.818682
R2126 iovss.n6 iovss.n5 0.818682
R2127 iovss.n217 iovss.n216 0.818682
R2128 iovss.n3 iovss.n2 0.818682
R2129 iovss.n85 iovss.n84 0.416993
R2130 iovss.n219 iovss.n218 0.416993
R2131 iovss.n90 iovss.n80 0.201704
R2132 iovss.n221 iovss.n220 0.2005
R2133 iovss.n215 iovss.n1 0.2005
R2134 iovss.n214 iovss.n213 0.2005
R2135 iovss.n11 iovss.n7 0.2005
R2136 iovss.n209 iovss.n208 0.2005
R2137 iovss.n200 iovss.n9 0.2005
R2138 iovss.n199 iovss.n198 0.2005
R2139 iovss.n20 iovss.n16 0.2005
R2140 iovss.n194 iovss.n193 0.2005
R2141 iovss.n185 iovss.n18 0.2005
R2142 iovss.n184 iovss.n183 0.2005
R2143 iovss.n29 iovss.n25 0.2005
R2144 iovss.n179 iovss.n178 0.2005
R2145 iovss.n170 iovss.n27 0.2005
R2146 iovss.n169 iovss.n168 0.2005
R2147 iovss.n38 iovss.n34 0.2005
R2148 iovss.n164 iovss.n163 0.2005
R2149 iovss.n155 iovss.n36 0.2005
R2150 iovss.n154 iovss.n153 0.2005
R2151 iovss.n47 iovss.n43 0.2005
R2152 iovss.n149 iovss.n148 0.2005
R2153 iovss.n140 iovss.n45 0.2005
R2154 iovss.n139 iovss.n138 0.2005
R2155 iovss.n56 iovss.n52 0.2005
R2156 iovss.n134 iovss.n133 0.2005
R2157 iovss.n125 iovss.n54 0.2005
R2158 iovss.n124 iovss.n123 0.2005
R2159 iovss.n65 iovss.n61 0.2005
R2160 iovss.n119 iovss.n118 0.2005
R2161 iovss.n110 iovss.n63 0.2005
R2162 iovss.n109 iovss.n108 0.2005
R2163 iovss.n74 iovss.n70 0.2005
R2164 iovss.n104 iovss.n103 0.2005
R2165 iovss.n95 iovss.n72 0.2005
R2166 iovss.n94 iovss.n93 0.2005
R2167 iovss.n82 iovss.n79 0.2005
R2168 iovss.n89 iovss.n88 0.2005
R2169 iovss.n222 iovss.n221 0.1105
R2170 iovss.n1 iovss.n0 0.1105
R2171 iovss.n213 iovss.n212 0.1105
R2172 iovss.n211 iovss.n7 0.1105
R2173 iovss.n210 iovss.n209 0.1105
R2174 iovss.n9 iovss.n8 0.1105
R2175 iovss.n198 iovss.n197 0.1105
R2176 iovss.n196 iovss.n16 0.1105
R2177 iovss.n195 iovss.n194 0.1105
R2178 iovss.n18 iovss.n17 0.1105
R2179 iovss.n183 iovss.n182 0.1105
R2180 iovss.n181 iovss.n25 0.1105
R2181 iovss.n180 iovss.n179 0.1105
R2182 iovss.n27 iovss.n26 0.1105
R2183 iovss.n168 iovss.n167 0.1105
R2184 iovss.n166 iovss.n34 0.1105
R2185 iovss.n165 iovss.n164 0.1105
R2186 iovss.n36 iovss.n35 0.1105
R2187 iovss.n153 iovss.n152 0.1105
R2188 iovss.n151 iovss.n43 0.1105
R2189 iovss.n150 iovss.n149 0.1105
R2190 iovss.n45 iovss.n44 0.1105
R2191 iovss.n138 iovss.n137 0.1105
R2192 iovss.n136 iovss.n52 0.1105
R2193 iovss.n135 iovss.n134 0.1105
R2194 iovss.n54 iovss.n53 0.1105
R2195 iovss.n123 iovss.n122 0.1105
R2196 iovss.n121 iovss.n61 0.1105
R2197 iovss.n120 iovss.n119 0.1105
R2198 iovss.n63 iovss.n62 0.1105
R2199 iovss.n108 iovss.n107 0.1105
R2200 iovss.n106 iovss.n70 0.1105
R2201 iovss.n105 iovss.n104 0.1105
R2202 iovss.n72 iovss.n71 0.1105
R2203 iovss.n93 iovss.n92 0.1105
R2204 iovss.n91 iovss.n79 0.1105
R2205 iovss.n91 iovss.n90 0.0568704
R2206 iovss.n85 iovss.n76 0.00740196
R2207 iovss.n98 iovss.n76 0.00740196
R2208 iovss.n99 iovss.n98 0.00740196
R2209 iovss.n100 iovss.n99 0.00740196
R2210 iovss.n100 iovss.n67 0.00740196
R2211 iovss.n113 iovss.n67 0.00740196
R2212 iovss.n114 iovss.n113 0.00740196
R2213 iovss.n115 iovss.n114 0.00740196
R2214 iovss.n115 iovss.n58 0.00740196
R2215 iovss.n128 iovss.n58 0.00740196
R2216 iovss.n129 iovss.n128 0.00740196
R2217 iovss.n130 iovss.n129 0.00740196
R2218 iovss.n130 iovss.n49 0.00740196
R2219 iovss.n143 iovss.n49 0.00740196
R2220 iovss.n144 iovss.n143 0.00740196
R2221 iovss.n145 iovss.n144 0.00740196
R2222 iovss.n145 iovss.n40 0.00740196
R2223 iovss.n158 iovss.n40 0.00740196
R2224 iovss.n159 iovss.n158 0.00740196
R2225 iovss.n160 iovss.n159 0.00740196
R2226 iovss.n160 iovss.n31 0.00740196
R2227 iovss.n173 iovss.n31 0.00740196
R2228 iovss.n174 iovss.n173 0.00740196
R2229 iovss.n175 iovss.n174 0.00740196
R2230 iovss.n175 iovss.n22 0.00740196
R2231 iovss.n188 iovss.n22 0.00740196
R2232 iovss.n189 iovss.n188 0.00740196
R2233 iovss.n190 iovss.n189 0.00740196
R2234 iovss.n190 iovss.n13 0.00740196
R2235 iovss.n203 iovss.n13 0.00740196
R2236 iovss.n204 iovss.n203 0.00740196
R2237 iovss.n205 iovss.n204 0.00740196
R2238 iovss.n205 iovss.n4 0.00740196
R2239 iovss.n218 iovss.n4 0.00740196
R2240 iovss.n86 iovss.n83 0.00740196
R2241 iovss.n86 iovss.n77 0.00740196
R2242 iovss.n97 iovss.n77 0.00740196
R2243 iovss.n97 iovss.n75 0.00740196
R2244 iovss.n101 iovss.n75 0.00740196
R2245 iovss.n101 iovss.n68 0.00740196
R2246 iovss.n112 iovss.n68 0.00740196
R2247 iovss.n112 iovss.n66 0.00740196
R2248 iovss.n116 iovss.n66 0.00740196
R2249 iovss.n116 iovss.n59 0.00740196
R2250 iovss.n127 iovss.n59 0.00740196
R2251 iovss.n127 iovss.n57 0.00740196
R2252 iovss.n131 iovss.n57 0.00740196
R2253 iovss.n131 iovss.n50 0.00740196
R2254 iovss.n142 iovss.n50 0.00740196
R2255 iovss.n142 iovss.n48 0.00740196
R2256 iovss.n146 iovss.n48 0.00740196
R2257 iovss.n146 iovss.n41 0.00740196
R2258 iovss.n157 iovss.n41 0.00740196
R2259 iovss.n157 iovss.n39 0.00740196
R2260 iovss.n161 iovss.n39 0.00740196
R2261 iovss.n161 iovss.n32 0.00740196
R2262 iovss.n172 iovss.n32 0.00740196
R2263 iovss.n172 iovss.n30 0.00740196
R2264 iovss.n176 iovss.n30 0.00740196
R2265 iovss.n176 iovss.n23 0.00740196
R2266 iovss.n187 iovss.n23 0.00740196
R2267 iovss.n187 iovss.n21 0.00740196
R2268 iovss.n191 iovss.n21 0.00740196
R2269 iovss.n191 iovss.n14 0.00740196
R2270 iovss.n202 iovss.n14 0.00740196
R2271 iovss.n202 iovss.n12 0.00740196
R2272 iovss.n206 iovss.n12 0.00740196
R2273 iovss.n206 iovss.n5 0.00740196
R2274 iovss.n217 iovss.n5 0.00740196
R2275 iovss.n217 iovss.n3 0.00740196
R2276 iovss.n219 iovss.n3 0.00442211
R2277 iovss.n84 iovss.n83 0.00442211
R2278 iovss.n81 iovss.n80 0.00395098
R2279 iovss.n88 iovss.n81 0.00395098
R2280 iovss.n88 iovss.n87 0.00395098
R2281 iovss.n87 iovss.n82 0.00395098
R2282 iovss.n82 iovss.n78 0.00395098
R2283 iovss.n94 iovss.n78 0.00395098
R2284 iovss.n96 iovss.n94 0.00395098
R2285 iovss.n96 iovss.n95 0.00395098
R2286 iovss.n95 iovss.n73 0.00395098
R2287 iovss.n103 iovss.n73 0.00395098
R2288 iovss.n103 iovss.n102 0.00395098
R2289 iovss.n102 iovss.n74 0.00395098
R2290 iovss.n74 iovss.n69 0.00395098
R2291 iovss.n109 iovss.n69 0.00395098
R2292 iovss.n111 iovss.n109 0.00395098
R2293 iovss.n111 iovss.n110 0.00395098
R2294 iovss.n110 iovss.n64 0.00395098
R2295 iovss.n118 iovss.n64 0.00395098
R2296 iovss.n118 iovss.n117 0.00395098
R2297 iovss.n117 iovss.n65 0.00395098
R2298 iovss.n65 iovss.n60 0.00395098
R2299 iovss.n124 iovss.n60 0.00395098
R2300 iovss.n126 iovss.n124 0.00395098
R2301 iovss.n126 iovss.n125 0.00395098
R2302 iovss.n125 iovss.n55 0.00395098
R2303 iovss.n133 iovss.n55 0.00395098
R2304 iovss.n133 iovss.n132 0.00395098
R2305 iovss.n132 iovss.n56 0.00395098
R2306 iovss.n56 iovss.n51 0.00395098
R2307 iovss.n139 iovss.n51 0.00395098
R2308 iovss.n141 iovss.n139 0.00395098
R2309 iovss.n141 iovss.n140 0.00395098
R2310 iovss.n140 iovss.n46 0.00395098
R2311 iovss.n148 iovss.n46 0.00395098
R2312 iovss.n148 iovss.n147 0.00395098
R2313 iovss.n147 iovss.n47 0.00395098
R2314 iovss.n47 iovss.n42 0.00395098
R2315 iovss.n154 iovss.n42 0.00395098
R2316 iovss.n156 iovss.n154 0.00395098
R2317 iovss.n156 iovss.n155 0.00395098
R2318 iovss.n155 iovss.n37 0.00395098
R2319 iovss.n163 iovss.n37 0.00395098
R2320 iovss.n163 iovss.n162 0.00395098
R2321 iovss.n162 iovss.n38 0.00395098
R2322 iovss.n38 iovss.n33 0.00395098
R2323 iovss.n169 iovss.n33 0.00395098
R2324 iovss.n171 iovss.n169 0.00395098
R2325 iovss.n171 iovss.n170 0.00395098
R2326 iovss.n170 iovss.n28 0.00395098
R2327 iovss.n178 iovss.n28 0.00395098
R2328 iovss.n178 iovss.n177 0.00395098
R2329 iovss.n177 iovss.n29 0.00395098
R2330 iovss.n29 iovss.n24 0.00395098
R2331 iovss.n184 iovss.n24 0.00395098
R2332 iovss.n186 iovss.n184 0.00395098
R2333 iovss.n186 iovss.n185 0.00395098
R2334 iovss.n185 iovss.n19 0.00395098
R2335 iovss.n193 iovss.n19 0.00395098
R2336 iovss.n193 iovss.n192 0.00395098
R2337 iovss.n192 iovss.n20 0.00395098
R2338 iovss.n20 iovss.n15 0.00395098
R2339 iovss.n199 iovss.n15 0.00395098
R2340 iovss.n201 iovss.n199 0.00395098
R2341 iovss.n201 iovss.n200 0.00395098
R2342 iovss.n200 iovss.n10 0.00395098
R2343 iovss.n208 iovss.n10 0.00395098
R2344 iovss.n208 iovss.n207 0.00395098
R2345 iovss.n207 iovss.n11 0.00395098
R2346 iovss.n11 iovss.n6 0.00395098
R2347 iovss.n214 iovss.n6 0.00395098
R2348 iovss.n216 iovss.n214 0.00395098
R2349 iovss.n216 iovss.n215 0.00395098
R2350 iovss.n215 iovss.n2 0.00395098
R2351 iovss.n220 iovss.n2 0.00395098
R2352 iovss.n221 iovss 0.00261765
R2353 iovss iovss.n222 0.00196667
R2354 iovss.n89 iovss.n79 0.00191176
R2355 iovss.n93 iovss.n79 0.00191176
R2356 iovss.n93 iovss.n72 0.00191176
R2357 iovss.n104 iovss.n72 0.00191176
R2358 iovss.n104 iovss.n70 0.00191176
R2359 iovss.n108 iovss.n70 0.00191176
R2360 iovss.n108 iovss.n63 0.00191176
R2361 iovss.n119 iovss.n63 0.00191176
R2362 iovss.n119 iovss.n61 0.00191176
R2363 iovss.n123 iovss.n61 0.00191176
R2364 iovss.n123 iovss.n54 0.00191176
R2365 iovss.n134 iovss.n54 0.00191176
R2366 iovss.n134 iovss.n52 0.00191176
R2367 iovss.n138 iovss.n52 0.00191176
R2368 iovss.n138 iovss.n45 0.00191176
R2369 iovss.n149 iovss.n45 0.00191176
R2370 iovss.n149 iovss.n43 0.00191176
R2371 iovss.n153 iovss.n43 0.00191176
R2372 iovss.n153 iovss.n36 0.00191176
R2373 iovss.n164 iovss.n36 0.00191176
R2374 iovss.n164 iovss.n34 0.00191176
R2375 iovss.n168 iovss.n34 0.00191176
R2376 iovss.n168 iovss.n27 0.00191176
R2377 iovss.n179 iovss.n27 0.00191176
R2378 iovss.n179 iovss.n25 0.00191176
R2379 iovss.n183 iovss.n25 0.00191176
R2380 iovss.n183 iovss.n18 0.00191176
R2381 iovss.n194 iovss.n18 0.00191176
R2382 iovss.n194 iovss.n16 0.00191176
R2383 iovss.n198 iovss.n16 0.00191176
R2384 iovss.n198 iovss.n9 0.00191176
R2385 iovss.n209 iovss.n9 0.00191176
R2386 iovss.n209 iovss.n7 0.00191176
R2387 iovss.n213 iovss.n7 0.00191176
R2388 iovss.n213 iovss.n1 0.00191176
R2389 iovss.n221 iovss.n1 0.00191176
R2390 iovss.n90 iovss.n89 0.0016983
R2391 iovss.n92 iovss.n91 0.00147778
R2392 iovss.n92 iovss.n71 0.00147778
R2393 iovss.n105 iovss.n71 0.00147778
R2394 iovss.n106 iovss.n105 0.00147778
R2395 iovss.n107 iovss.n106 0.00147778
R2396 iovss.n107 iovss.n62 0.00147778
R2397 iovss.n120 iovss.n62 0.00147778
R2398 iovss.n121 iovss.n120 0.00147778
R2399 iovss.n122 iovss.n121 0.00147778
R2400 iovss.n122 iovss.n53 0.00147778
R2401 iovss.n135 iovss.n53 0.00147778
R2402 iovss.n136 iovss.n135 0.00147778
R2403 iovss.n137 iovss.n136 0.00147778
R2404 iovss.n137 iovss.n44 0.00147778
R2405 iovss.n150 iovss.n44 0.00147778
R2406 iovss.n151 iovss.n150 0.00147778
R2407 iovss.n152 iovss.n151 0.00147778
R2408 iovss.n152 iovss.n35 0.00147778
R2409 iovss.n165 iovss.n35 0.00147778
R2410 iovss.n166 iovss.n165 0.00147778
R2411 iovss.n167 iovss.n166 0.00147778
R2412 iovss.n167 iovss.n26 0.00147778
R2413 iovss.n180 iovss.n26 0.00147778
R2414 iovss.n181 iovss.n180 0.00147778
R2415 iovss.n182 iovss.n181 0.00147778
R2416 iovss.n182 iovss.n17 0.00147778
R2417 iovss.n195 iovss.n17 0.00147778
R2418 iovss.n196 iovss.n195 0.00147778
R2419 iovss.n197 iovss.n196 0.00147778
R2420 iovss.n197 iovss.n8 0.00147778
R2421 iovss.n210 iovss.n8 0.00147778
R2422 iovss.n211 iovss.n210 0.00147778
R2423 iovss.n212 iovss.n211 0.00147778
R2424 iovss.n212 iovss.n0 0.00147778
R2425 iovss.n222 iovss.n0 0.00147778
R2426 c2p_en.n2 c2p_en.t0 15.0005
R2427 c2p_en.n1 c2p_en.t1 15.0005
R2428 c2p_en.n4 c2p_en.n1 9.74312
R2429 c2p_en.n3 c2p_en.n2 9.22574
R2430 c2p_en.n0 c2p_en 9.10188
R2431 c2p_en.n2 c2p_en 2.16907
R2432 c2p_en.n1 c2p_en 2.16907
R2433 c2p_en.n4 c2p_en.n0 1.63153
R2434 c2p_en.n0 c2p_en 0.99754
R2435 c2p_en c2p_en.n4 0.0885
R2436 c2p_en.n3 c2p_en 0.0308448
R2437 c2p_en.n4 c2p_en.n3 0.0141552
R2438 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t3 21.2194
R2439 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n0 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t2 15.755
R2440 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n1 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n0 12.6797
R2441 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n0 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq 1.8683
R2442 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n3 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t0 1.73646
R2443 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n3 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n2 1.57533
R2444 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n2 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t1 1.43953
R2445 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n2 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n1 0.782552
R2446 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n3 0.753577
R2447 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n1 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq 0.0764524
R2448 c2p.n2 c2p.t1 15.0005
R2449 c2p.n1 c2p.t0 15.0005
R2450 c2p.n4 c2p.n1 12.0592
R2451 c2p.n3 c2p.n2 11.3445
R2452 c2p.n0 c2p 9.10188
R2453 c2p.n2 c2p 2.16907
R2454 c2p.n1 c2p 2.16907
R2455 c2p.n4 c2p.n0 0.404086
R2456 c2p.n0 c2p 0.28562
R2457 c2p c2p.n4 0.0885
R2458 c2p.n3 c2p 0.0308448
R2459 c2p.n4 c2p.n3 0.0141552
C0 vdd a_4358_31526# 0.81747f
C1 vdd c2p 1.52081f
C2 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq a_4358_31526# 0.99584f
C3 sg13g2_DCNDiode_0.guard pad 7.46684f
C4 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq c2p 0.43902f
C5 iovdd sg13g2_LevelDown_0.sg13g2_SecondaryProtection_0.core 1.37355f
C6 vdd p2c 2.6001f
C7 vdd sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq 2.11533f
C8 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq a_4426_30170# 0.1286f
C9 a_12038_31490# sg13g2_LevelDown_0.sg13g2_SecondaryProtection_0.core 0.31408f
C10 a_3724_30170# iovdd 0.84924f
C11 iovdd a_4358_30206# 0.28407f
C12 vdd sg13g2_LevelDown_0.sg13g2_SecondaryProtection_0.core 0.51442f
C13 a_3724_30170# sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq 0.1286f
C14 p2c sg13g2_LevelDown_0.sg13g2_SecondaryProtection_0.core 0.10336f
C15 c2p_en sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq 1.6012f
C16 a_4358_31526# a_4358_30206# 0.15491f
C17 sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq 1.30685f
C18 c2p c2p_en 0.53273f
C19 sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq a_3656_31526# 0.99218f
C20 a_3656_30206# iovdd 0.30461f
C21 vdd c2p_en 1.46533f
C22 iovdd a_4426_30170# 0.84126f
C23 a_3724_30170# a_3656_30206# 0.37106f
C24 sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq a_4358_31526# 0.30586f
C25 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq c2p_en 1.59673f
C26 sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq c2p 0.65338f
C27 a_4358_30206# a_4426_30170# 0.37106f
C28 a_12038_31490# vdd 1.10866f
C29 vdd sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq 1.87035f
C30 c2p sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq 0.56766f
C31 iovdd pad 47.63779f
C32 a_12038_31490# p2c 0.25311f
C33 vdd sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq 1.00261f
C34 vdd a_3656_31526# 0.79605f
C35 a_3656_30206# a_3656_31526# 0.15491f
C36 pad iovss 0.13534p
C37 p2c iovss 1.03179f
C38 c2p_en iovss 2.18641f
C39 c2p iovss 2.43746f
C40 iovdd iovss 0.14274p
C41 vdd iovss 0.24597p
C42 a_12137_28308# iovss 0.47362f $ **FLOATING
C43 a_4358_30206# iovss 0.23648f
C44 a_3656_30206# iovss 0.45339f
C45 a_4426_30170# iovss 1.28302f
C46 a_3724_30170# iovss 1.27692f
C47 sg13g2_LevelDown_0.sg13g2_SecondaryProtection_0.core iovss 6.27806f
C48 a_4358_31526# iovss 1.33907f
C49 a_3656_31526# iovss 1.89714f
C50 a_12038_31490# iovss 1.36953f
C51 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq iovss 2.98668f
C52 sg13g2_GateDecode_0.sg13g2_io_nor2_x1_0.nq iovss 2.73965f
C53 sg13g2_GateDecode_0.sg13g2_io_inv_x1_0.nq iovss 1.32815f
C54 sg13g2_DCNDiode_0.guard iovss 53.69175f $ **FLOATING
C55 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t1 iovss 0.16985f
C56 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t3 iovss 0.12361f
C57 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t2 iovss 0.16083f
C58 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n0 iovss 0.78384f
C59 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.t0 iovss 0.23765f
C60 sg13g2_GateDecode_0.sg13g2_io_nand2_x1_0.nq.n3 iovss 0.5473f
C61 sg13g2_GateDecode_0.ngate.t0 iovss 0.11359f
C62 sg13g2_GateDecode_0.ngate.t1 iovss 0.22122f
C63 sg13g2_GateDecode_0.ngate.n0 iovss 0.26675f
C64 sg13g2_Clamp_N15N15D_0.gate iovss 3.7933f
C65 sg13g2_GateDecode_0.ngate.t3 iovss 0.47567f
C66 sg13g2_GateDecode_0.ngate.t15 iovss 0.46415f
C67 sg13g2_GateDecode_0.ngate.n1 iovss 0.2535f
C68 sg13g2_GateDecode_0.ngate.t11 iovss 0.46415f
C69 sg13g2_GateDecode_0.ngate.n2 iovss 0.14203f
C70 sg13g2_GateDecode_0.ngate.t5 iovss 0.46415f
C71 sg13g2_GateDecode_0.ngate.n3 iovss 0.14203f
C72 sg13g2_GateDecode_0.ngate.t9 iovss 0.46415f
C73 sg13g2_GateDecode_0.ngate.n4 iovss 0.14203f
C74 sg13g2_GateDecode_0.ngate.t8 iovss 0.46415f
C75 sg13g2_GateDecode_0.ngate.n5 iovss 0.14203f
C76 sg13g2_GateDecode_0.ngate.t16 iovss 0.46415f
C77 sg13g2_GateDecode_0.ngate.n6 iovss 0.14203f
C78 sg13g2_GateDecode_0.ngate.t6 iovss 0.46415f
C79 sg13g2_GateDecode_0.ngate.n7 iovss 0.14203f
C80 sg13g2_GateDecode_0.ngate.t17 iovss 0.46415f
C81 sg13g2_GateDecode_0.ngate.n8 iovss 0.14203f
C82 sg13g2_GateDecode_0.ngate.t14 iovss 0.46415f
C83 sg13g2_GateDecode_0.ngate.n9 iovss 0.14203f
C84 sg13g2_GateDecode_0.ngate.t4 iovss 0.46415f
C85 sg13g2_GateDecode_0.ngate.n10 iovss 0.14203f
C86 sg13g2_GateDecode_0.ngate.t13 iovss 0.46415f
C87 sg13g2_GateDecode_0.ngate.n11 iovss 0.14203f
C88 sg13g2_GateDecode_0.ngate.t7 iovss 0.46415f
C89 sg13g2_GateDecode_0.ngate.n12 iovss 0.14203f
C90 sg13g2_GateDecode_0.ngate.t2 iovss 0.46415f
C91 sg13g2_GateDecode_0.ngate.n13 iovss 0.14203f
C92 sg13g2_GateDecode_0.ngate.t10 iovss 0.46415f
C93 sg13g2_GateDecode_0.ngate.n14 iovss 0.29439f
C94 sg13g2_GateDecode_0.ngate.n15 iovss 0.22009f
C95 sg13g2_GateDecode_0.sg13g2_LevelUp_0.o iovss 2.72464f
C96 pad.t4 iovss 0.20893f
C97 pad.n0 iovss 0.19654f
C98 pad.n28 iovss 0.21184f
C99 pad.n29 iovss 0.21184f
C100 pad.n30 iovss 0.21184f
C101 pad.n31 iovss 0.21184f
C102 pad.n32 iovss 0.21184f
C103 pad.n33 iovss 0.21184f
C104 pad.n34 iovss 0.21184f
C105 pad.n35 iovss 0.21184f
C106 pad.n36 iovss 0.21184f
C107 pad.n37 iovss 0.21184f
C108 pad.n38 iovss 0.21184f
C109 pad.n39 iovss 0.21184f
C110 pad.n40 iovss 0.21184f
C111 pad.n41 iovss 0.21184f
C112 pad.n42 iovss 0.21184f
C113 pad.n43 iovss 0.21184f
C114 pad.n44 iovss 0.21184f
C115 pad.n45 iovss 0.21184f
C116 pad.n46 iovss 0.21184f
C117 pad.n47 iovss 0.21184f
C118 pad.n48 iovss 0.21184f
C119 pad.n49 iovss 0.21184f
C120 pad.n53 iovss 0.38251f
C121 pad.n55 iovss 0.10467f
C122 pad.n56 iovss 0.17875f
C123 pad.n62 iovss 0.38251f
C124 pad.n79 iovss 0.21184f
C125 pad.n80 iovss 0.21184f
C126 pad.n81 iovss 0.21184f
C127 pad.n82 iovss 0.21184f
C128 pad.n83 iovss 0.21184f
C129 pad.n84 iovss 0.21184f
C130 pad.n85 iovss 0.21184f
C131 pad.n86 iovss 0.21184f
C132 pad.n87 iovss 0.21184f
C133 pad.n88 iovss 0.21184f
C134 pad.n89 iovss 0.21184f
C135 pad.n90 iovss 0.21184f
C136 pad.n91 iovss 0.21184f
C137 pad.n92 iovss 0.21184f
C138 pad.n93 iovss 0.21184f
C139 pad.n94 iovss 0.21184f
C140 pad.n103 iovss 0.21184f
C141 pad.n104 iovss 0.21184f
C142 pad.n105 iovss 0.21184f
C143 pad.n106 iovss 0.21184f
C144 pad.n107 iovss 0.21184f
C145 pad.n108 iovss 0.21184f
C146 pad.n109 iovss 0.21184f
C147 pad.n118 iovss 0.21184f
C148 pad.n119 iovss 0.21184f
C149 pad.n120 iovss 0.21184f
C150 pad.n121 iovss 0.62857f
C151 pad.n122 iovss 0.21184f
C152 pad.n123 iovss 0.21184f
C153 pad.n124 iovss 0.21184f
C154 pad.n131 iovss 0.2127f
C155 pad.n132 iovss 0.21247f
C156 pad.n133 iovss 0.21818f
C157 pad.n134 iovss 0.21184f
C158 pad.n135 iovss 0.21184f
C159 pad.n136 iovss 0.21184f
C160 pad.n138 iovss 0.26586f
C161 pad.n139 iovss 0.32206f
C162 pad.n166 iovss 0.21184f
C163 pad.n167 iovss 0.21184f
C164 pad.n168 iovss 0.21184f
C165 pad.n169 iovss 0.21184f
C166 pad.n170 iovss 0.21184f
C167 pad.n171 iovss 0.21184f
C168 pad.n172 iovss 0.21184f
C169 pad.n173 iovss 0.21184f
C170 pad.n174 iovss 0.21184f
C171 pad.n203 iovss 0.21184f
C172 pad.n204 iovss 0.21184f
C173 pad.n205 iovss 0.21184f
C174 pad.n206 iovss 0.21184f
C175 pad.n207 iovss 0.21184f
C176 pad.n208 iovss 0.21184f
C177 pad.n209 iovss 0.21184f
C178 pad.n210 iovss 0.21184f
C179 pad.n211 iovss 0.21184f
C180 pad.n227 iovss 0.3859f
C181 pad.t25 iovss 1.24564f
C182 pad.t7 iovss 0.45548f
C183 pad.t9 iovss 0.32056f
C184 pad.n229 iovss 0.37719f
C185 pad.n230 iovss 0.13036f
C186 pad.n233 iovss 0.17875f
C187 pad.t16 iovss 0.45548f
C188 pad.t18 iovss 0.32056f
C189 pad.n238 iovss 0.37719f
C190 pad.n239 iovss 0.13036f
C191 pad.n241 iovss 0.15065f
C192 pad.t17 iovss 0.45548f
C193 pad.t8 iovss 0.32056f
C194 pad.n244 iovss 0.37719f
C195 pad.t19 iovss 0.45548f
C196 pad.t20 iovss 0.32056f
C197 pad.n246 iovss 0.37719f
C198 pad.n248 iovss 0.38251f
C199 pad.n249 iovss 0.13036f
C200 pad.t21 iovss 0.21709f
C201 pad.n251 iovss 1.01081f
C202 pad.t22 iovss 0.21709f
C203 pad.n252 iovss 0.20682f
C204 pad.n253 iovss 0.13375f
C205 pad.n254 iovss 0.17875f
C206 pad.t11 iovss 0.45548f
C207 pad.t12 iovss 0.32056f
C208 pad.n257 iovss 0.37719f
C209 pad.n258 iovss 0.15065f
C210 pad.n262 iovss 0.10467f
C211 pad.n263 iovss 0.38251f
C212 pad.n264 iovss 0.10467f
C213 pad.n265 iovss 0.38251f
C214 pad.n266 iovss 0.13036f
C215 pad.n267 iovss 0.10467f
C216 pad.t14 iovss 0.45548f
C217 pad.t15 iovss 0.32056f
C218 pad.n270 iovss 0.37719f
C219 pad.t3 iovss 0.20893f
C220 pad.n271 iovss 0.19654f
C221 pad.n273 iovss 0.15065f
C222 pad.n275 iovss 0.38251f
C223 pad.n276 iovss 0.38251f
C224 pad.n277 iovss 0.13036f
C225 pad.t10 iovss 0.45548f
C226 pad.t13 iovss 0.32056f
C227 pad.n281 iovss 0.37719f
C228 pad.n282 iovss 0.10131f
C229 pad.n283 iovss 0.38251f
C230 pad.n284 iovss 0.13036f
C231 pad.n285 iovss 0.10131f
C232 pad.t27 iovss 1.24564f
C233 pad.n289 iovss 0.13036f
C234 pad.n291 iovss 0.38251f
C235 pad.t23 iovss 0.20893f
C236 pad.n296 iovss 0.19654f
C237 pad.t6 iovss 0.20893f
C238 pad.n317 iovss 0.19654f
C239 pad.n319 iovss 0.15065f
C240 pad.n320 iovss 0.38251f
C241 pad.n324 iovss 0.38251f
C242 pad.n325 iovss 0.38251f
C243 pad.t26 iovss 1.24564f
C244 pad.n330 iovss 0.38251f
C245 pad.t5 iovss 0.20893f
C246 pad.n331 iovss 0.19654f
C247 pad.n332 iovss 0.15065f
C248 pad.n333 iovss 0.38251f
C249 pad.n336 iovss 0.10131f
C250 pad.n337 iovss 0.17875f
C251 pad.n338 iovss 0.3859f
C252 pad.n339 iovss 0.15405f
C253 pad.t2 iovss 0.14057f
C254 pad.n340 iovss 0.19654f
C255 pad.n358 iovss 0.21184f
C256 pad.n359 iovss 0.21184f
C257 pad.n360 iovss 0.21184f
C258 pad.n361 iovss 0.21184f
C259 pad.n362 iovss 0.21184f
C260 pad.n363 iovss 0.21184f
C261 pad.n364 iovss 0.21184f
C262 pad.n365 iovss 0.21184f
C263 pad.n366 iovss 0.21184f
C264 pad.n367 iovss 0.21184f
C265 pad.n368 iovss 0.21184f
C266 pad.n369 iovss 0.21184f
C267 pad.n370 iovss 0.21184f
C268 pad.n371 iovss 0.21184f
C269 pad.n372 iovss 0.21184f
C270 pad.n373 iovss 0.21184f
C271 pad.n374 iovss 0.21184f
C272 pad.n375 iovss 0.21184f
C273 pad.n376 iovss 0.21184f
C274 pad.n377 iovss 0.21184f
C275 pad.t1 iovss 0.20893f
C276 pad.n406 iovss 0.19654f
C277 pad.n407 iovss 0.15065f
C278 pad.n408 iovss 0.10131f
C279 pad.t28 iovss 1.24564f
C280 pad.n412 iovss 0.15065f
C281 pad.t0 iovss 0.20893f
C282 pad.n413 iovss 0.19654f
C283 pad.n431 iovss 0.21184f
C284 pad.n432 iovss 0.21184f
C285 pad.n433 iovss 0.21184f
C286 pad.n434 iovss 0.21184f
C287 pad.n435 iovss 0.21184f
C288 pad.n436 iovss 0.21184f
C289 pad.n437 iovss 0.21184f
C290 pad.n438 iovss 0.21184f
C291 pad.n439 iovss 0.21184f
C292 pad.n440 iovss 0.21184f
C293 pad.n441 iovss 0.21184f
C294 pad.n442 iovss 0.21184f
C295 pad.n443 iovss 0.21184f
C296 pad.n444 iovss 0.21184f
C297 pad.n445 iovss 0.21184f
C298 pad.n446 iovss 0.21184f
C299 pad.n447 iovss 0.21184f
C300 pad.n448 iovss 0.21184f
C301 pad.n449 iovss 0.21184f
C302 pad.n450 iovss 0.21184f
C303 pad.n451 iovss 0.21184f
C304 pad.n452 iovss 0.21184f
C305 pad.n453 iovss 0.21184f
C306 pad.n454 iovss 0.21184f
C307 pad.n455 iovss 0.21184f
C308 pad.n456 iovss 0.21184f
C309 pad.n457 iovss 0.21184f
C310 pad.n458 iovss 0.21184f
C311 pad.n459 iovss 0.21184f
C312 pad.n460 iovss 0.32207f
C313 pad.n477 iovss 0.21184f
C314 pad.n486 iovss 0.26584f
C315 pad.n487 iovss 0.2127f
C316 pad.n488 iovss 0.21184f
C317 pad.n489 iovss 0.15888f
C318 pad.n490 iovss 0.21184f
C319 pad.n491 iovss 0.21184f
C320 pad.n492 iovss 0.21184f
C321 pad.n493 iovss 0.21184f
C322 pad.n494 iovss 0.21184f
C323 pad.n495 iovss 0.21184f
C324 pad.n496 iovss 0.21184f
C325 pad.n497 iovss 0.21184f
C326 pad.n498 iovss 0.21184f
C327 iovdd.t14 iovss 10.7651f
C328 iovdd.n75 iovss 0.50981f
C329 iovdd.n121 iovss 0.31591f
C330 iovdd.n122 iovss 0.41842f
C331 iovdd.n123 iovss 0.41842f
C332 iovdd.n124 iovss 0.41842f
C333 iovdd.n125 iovss 0.20921f
C334 iovdd.n126 iovss 0.20921f
C335 iovdd.n127 iovss 0.41842f
C336 iovdd.n128 iovss 0.3692f
C337 iovdd.n129 iovss 0.41842f
C338 iovdd.n130 iovss 0.20921f
C339 iovdd.n131 iovss 0.41842f
C340 iovdd.n132 iovss 0.284f
C341 iovdd.n134 iovss 0.20766f
C342 iovdd.n135 iovss 0.41842f
C343 iovdd.n136 iovss 0.20921f
C344 iovdd.n137 iovss 0.20921f
C345 iovdd.n138 iovss 0.41842f
C346 iovdd.n139 iovss 0.3692f
C347 iovdd.n140 iovss 0.41842f
C348 iovdd.n141 iovss 0.20921f
C349 iovdd.n142 iovss 0.41842f
C350 iovdd.n143 iovss 0.31591f
C351 iovdd.n145 iovss 0.29237f
C352 iovdd.n146 iovss 0.41842f
C353 iovdd.n147 iovss 0.20921f
C354 iovdd.n148 iovss 0.20921f
C355 iovdd.n149 iovss 0.41842f
C356 iovdd.n150 iovss 0.3692f
C357 iovdd.n151 iovss 0.41842f
C358 iovdd.n152 iovss 0.20921f
C359 iovdd.n153 iovss 0.41842f
C360 iovdd.n154 iovss 0.41842f
C361 iovdd.n155 iovss 0.41842f
C362 iovdd.n156 iovss 0.20921f
C363 iovdd.n157 iovss 0.20921f
C364 iovdd.n158 iovss 0.41842f
C365 iovdd.n159 iovss 0.3692f
C366 iovdd.n160 iovss 0.41842f
C367 iovdd.n161 iovss 0.20921f
C368 iovdd.n162 iovss 0.41842f
C369 iovdd.n163 iovss 0.41842f
C370 iovdd.n164 iovss 0.41842f
C371 iovdd.n165 iovss 0.20921f
C372 iovdd.n166 iovss 0.20921f
C373 iovdd.n167 iovss 0.41842f
C374 iovdd.n168 iovss 0.3692f
C375 iovdd.n169 iovss 0.41842f
C376 iovdd.n170 iovss 0.20921f
C377 iovdd.n171 iovss 0.41842f
C378 iovdd.n172 iovss 0.41842f
C379 iovdd.n173 iovss 0.41842f
C380 iovdd.n174 iovss 0.20921f
C381 iovdd.n175 iovss 0.20921f
C382 iovdd.n176 iovss 0.41842f
C383 iovdd.n177 iovss 1.45118f
C384 iovdd.n178 iovss 0.41842f
C385 iovdd.n179 iovss 0.20921f
C386 iovdd.n180 iovss 0.41842f
C387 iovdd.n181 iovss 0.73813f
C388 iovdd.n182 iovss 0.20921f
C389 iovdd.n183 iovss 0.8574f
C390 iovdd.n184 iovss 0.41842f
C391 iovdd.n185 iovss 0.20921f
C392 iovdd.n186 iovss 0.20921f
C393 iovdd.n187 iovss 0.41842f
C394 iovdd.n188 iovss 0.64929f
C395 iovdd.n189 iovss 1.44198f
C396 iovdd.n190 iovss 0.41842f
C397 iovdd.n191 iovss 0.41842f
C398 iovdd.n192 iovss 0.20921f
C399 iovdd.n193 iovss 0.20921f
C400 iovdd.n194 iovss 0.20921f
C401 iovdd.n195 iovss 0.41842f
C402 iovdd.n196 iovss 0.3692f
C403 iovdd.n197 iovss 0.3692f
C404 iovdd.n198 iovss 0.3692f
C405 iovdd.n199 iovss 0.41842f
C406 iovdd.n200 iovss 0.20921f
C407 iovdd.n201 iovss 0.20921f
C408 iovdd.n202 iovss 0.41842f
C409 iovdd.n203 iovss 0.41842f
C410 iovdd.n204 iovss 0.41842f
C411 iovdd.n205 iovss 0.41842f
C412 iovdd.n206 iovss 0.41842f
C413 iovdd.n207 iovss 0.20921f
C414 iovdd.n208 iovss 0.20921f
C415 iovdd.n209 iovss 0.20921f
C416 iovdd.n210 iovss 0.41842f
C417 iovdd.n211 iovss 0.3692f
C418 iovdd.n212 iovss 0.3692f
C419 iovdd.n213 iovss 0.3692f
C420 iovdd.n214 iovss 0.41842f
C421 iovdd.n215 iovss 0.20921f
C422 iovdd.n216 iovss 0.20921f
C423 iovdd.n217 iovss 0.41842f
C424 iovdd.n218 iovss 0.41842f
C425 iovdd.n219 iovss 0.41842f
C426 iovdd.n220 iovss 0.41842f
C427 iovdd.n221 iovss 0.41842f
C428 iovdd.n222 iovss 0.20921f
C429 iovdd.n223 iovss 0.20921f
C430 iovdd.n224 iovss 0.20921f
C431 iovdd.n225 iovss 0.41842f
C432 iovdd.n226 iovss 0.3692f
C433 iovdd.n227 iovss 0.3692f
C434 iovdd.n228 iovss 0.3692f
C435 iovdd.n229 iovss 0.41842f
C436 iovdd.n230 iovss 0.20921f
C437 iovdd.n231 iovss 0.20921f
C438 iovdd.n232 iovss 0.41842f
C439 iovdd.n233 iovss 0.41842f
C440 iovdd.n234 iovss 0.22856f
C441 iovdd.n235 iovss 0.20766f
C442 iovdd.n237 iovss 0.1751f
C443 iovdd.n246 iovss 0.20766f
C444 iovdd.n247 iovss 0.31591f
C445 iovdd.n248 iovss 0.41842f
C446 iovdd.n249 iovss 0.20921f
C447 iovdd.n250 iovss 0.20921f
C448 iovdd.n251 iovss 0.20921f
C449 iovdd.n252 iovss 0.41842f
C450 iovdd.n253 iovss 0.3692f
C451 iovdd.n254 iovss 0.3692f
C452 iovdd.n255 iovss 0.3692f
C453 iovdd.n256 iovss 0.41842f
C454 iovdd.n257 iovss 0.20921f
C455 iovdd.n258 iovss 0.20921f
C456 iovdd.n259 iovss 0.41842f
C457 iovdd.n260 iovss 0.23275f
C458 iovdd.n261 iovss 0.20766f
C459 iovdd.n280 iovss 0.20766f
C460 iovdd.n281 iovss 0.23693f
C461 iovdd.n282 iovss 0.28819f
C462 iovdd.n283 iovss 0.41842f
C463 iovdd.n284 iovss 0.20921f
C464 iovdd.n285 iovss 0.20921f
C465 iovdd.n286 iovss 0.20921f
C466 iovdd.n287 iovss 0.41842f
C467 iovdd.n288 iovss 0.3692f
C468 iovdd.n289 iovss 0.3692f
C469 iovdd.n290 iovss 0.3692f
C470 iovdd.n291 iovss 0.41842f
C471 iovdd.n292 iovss 0.20921f
C472 iovdd.n293 iovss 0.20921f
C473 iovdd.n294 iovss 0.41842f
C474 iovdd.n295 iovss 0.31591f
C475 iovdd.n296 iovss 0.20766f
C476 iovdd.n307 iovss 0.20766f
C477 iovdd.n308 iovss 0.24112f
C478 iovdd.n309 iovss 0.41842f
C479 iovdd.n310 iovss 0.20921f
C480 iovdd.n311 iovss 0.20921f
C481 iovdd.n312 iovss 0.20921f
C482 iovdd.n313 iovss 0.41842f
C483 iovdd.n314 iovss 0.3692f
C484 iovdd.n315 iovss 0.3692f
C485 iovdd.n316 iovss 0.3692f
C486 iovdd.n317 iovss 0.3692f
C487 iovdd.n318 iovss 0.41842f
C488 iovdd.n319 iovss 0.20921f
C489 iovdd.n320 iovss 0.41842f
C490 iovdd.n321 iovss 0.41842f
C491 iovdd.n322 iovss 0.41842f
C492 iovdd.n323 iovss 0.20921f
C493 iovdd.n324 iovss 0.3692f
C494 iovdd.n325 iovss 0.3692f
C495 iovdd.n326 iovss 0.3692f
C496 iovdd.n327 iovss 0.41842f
C497 iovdd.n328 iovss 0.20921f
C498 iovdd.n329 iovss 0.41842f
C499 iovdd.n330 iovss 0.41842f
C500 iovdd.n331 iovss 0.41842f
C501 iovdd.n332 iovss 0.41842f
C502 iovdd.n333 iovss 0.20921f
C503 iovdd.n334 iovss 0.3692f
C504 iovdd.n335 iovss 0.3692f
C505 iovdd.n336 iovss 0.3692f
C506 iovdd.n337 iovss 0.41842f
C507 iovdd.n338 iovss 0.20921f
C508 iovdd.n339 iovss 0.41842f
C509 iovdd.n340 iovss 0.41842f
C510 iovdd.n341 iovss 0.41842f
C511 iovdd.n342 iovss 0.41842f
C512 iovdd.n343 iovss 0.20921f
C513 iovdd.n344 iovss 0.3692f
C514 iovdd.n345 iovss 0.3692f
C515 iovdd.n346 iovss 0.3692f
C516 iovdd.n347 iovss 0.41842f
C517 iovdd.n348 iovss 0.20921f
C518 iovdd.n349 iovss 0.41842f
C519 iovdd.n350 iovss 1.44198f
C520 iovdd.n351 iovss 0.64929f
C521 iovdd.n352 iovss 0.3692f
C522 iovdd.n353 iovss 0.4615f
C523 iovdd.n354 iovss 0.52303f
C524 iovdd.n355 iovss 0.73308f
C525 iovdd.n356 iovss 0.20921f
C526 iovdd.n357 iovss 0.41842f
C527 iovdd.n358 iovss 0.41842f
C528 iovdd.n359 iovss 0.20921f
C529 iovdd.n360 iovss 0.20921f
C530 iovdd.n361 iovss 0.41842f
C531 iovdd.n362 iovss 0.41842f
C532 iovdd.n363 iovss 0.20921f
C533 iovdd.n364 iovss 0.20921f
C534 iovdd.n365 iovss 0.41842f
C535 iovdd.n366 iovss 0.41842f
C536 iovdd.n367 iovss 0.20921f
C537 iovdd.n368 iovss 0.20921f
C538 iovdd.n369 iovss 0.41842f
C539 iovdd.n370 iovss 0.41842f
C540 iovdd.n371 iovss 0.20921f
C541 iovdd.n372 iovss 0.20921f
C542 iovdd.n373 iovss 0.41842f
C543 iovdd.n374 iovss 0.41842f
C544 iovdd.n375 iovss 0.20921f
C545 iovdd.n376 iovss 0.20921f
C546 iovdd.n377 iovss 0.41842f
C547 iovdd.n378 iovss 0.41842f
C548 iovdd.n379 iovss 0.20921f
C549 iovdd.n380 iovss 0.20921f
C550 iovdd.n381 iovss 0.41842f
C551 iovdd.n382 iovss 0.41842f
C552 iovdd.n383 iovss 0.20921f
C553 iovdd.n384 iovss 0.20921f
C554 iovdd.n385 iovss 0.41842f
C555 iovdd.n386 iovss 0.41842f
C556 iovdd.n387 iovss 0.20921f
C557 iovdd.n388 iovss 0.20921f
C558 iovdd.n389 iovss 0.41842f
C559 iovdd.n390 iovss 0.27982f
C560 iovdd.n391 iovss 0.20766f
C561 iovdd.n398 iovss 0.12535f
C562 iovdd.n400 iovss 0.19586f
C563 iovdd.n422 iovss 0.12822f
C564 iovdd.t0 iovss 3.23621f
C565 iovdd.n511 iovss 0.83906f
C566 sg13g2_GateDecode_0.pgate.t0 iovss 0.25384f
C567 sg13g2_GateDecode_0.pgate.t1 iovss 0.49435f
C568 sg13g2_GateDecode_0.pgate.n0 iovss 0.59609f
C569 sg13g2_GateDecode_0.pgate.t5 iovss 3.09338f
C570 sg13g2_GateDecode_0.pgate.t16 iovss 3.09338f
C571 sg13g2_GateDecode_0.pgate.t10 iovss 3.09338f
C572 sg13g2_GateDecode_0.pgate.t4 iovss 3.09338f
C573 sg13g2_GateDecode_0.pgate.t11 iovss 3.09338f
C574 sg13g2_GateDecode_0.pgate.t3 iovss 3.09338f
C575 sg13g2_GateDecode_0.pgate.t12 iovss 3.09338f
C576 sg13g2_GateDecode_0.pgate.t8 iovss 3.09338f
C577 sg13g2_GateDecode_0.pgate.t14 iovss 3.09338f
C578 sg13g2_GateDecode_0.pgate.t6 iovss 3.09338f
C579 sg13g2_GateDecode_0.pgate.t17 iovss 3.09338f
C580 sg13g2_GateDecode_0.pgate.t9 iovss 3.09338f
C581 sg13g2_GateDecode_0.pgate.t15 iovss 3.09338f
C582 sg13g2_GateDecode_0.pgate.t13 iovss 3.09338f
C583 sg13g2_GateDecode_0.pgate.t7 iovss 3.1529f
C584 sg13g2_GateDecode_0.pgate.n2 iovss 1.09171f
C585 sg13g2_GateDecode_0.pgate.n3 iovss 0.59689f
C586 sg13g2_GateDecode_0.pgate.n4 iovss 0.59689f
C587 sg13g2_GateDecode_0.pgate.n5 iovss 0.59689f
C588 sg13g2_GateDecode_0.pgate.n6 iovss 0.59689f
C589 sg13g2_GateDecode_0.pgate.n7 iovss 0.59689f
C590 sg13g2_GateDecode_0.pgate.n8 iovss 0.59689f
C591 sg13g2_GateDecode_0.pgate.n9 iovss 0.59689f
C592 sg13g2_GateDecode_0.pgate.n10 iovss 0.59689f
C593 sg13g2_GateDecode_0.pgate.n11 iovss 0.59689f
C594 sg13g2_GateDecode_0.pgate.n12 iovss 0.59689f
C595 sg13g2_GateDecode_0.pgate.n13 iovss 0.59689f
C596 sg13g2_GateDecode_0.pgate.n14 iovss 0.59689f
C597 sg13g2_GateDecode_0.pgate.n15 iovss 0.93073f
C598 sg13g2_GateDecode_0.pgate.t2 iovss 0.20003f
C599 sg13g2_GateDecode_0.pgate.n16 iovss 0.10773f
C600 sg13g2_GateDecode_0.pgate.n17 iovss 0.38941f
C601 sg13g2_GateDecode_0.pgate.n18 iovss 2.90898f
C602 sg13g2_GateDecode_0.sg13g2_LevelUp_1.o iovss 2.67589f
C603 vdd.t0 iovss 0.16194f
C604 vdd.n41 iovss 0.13956f
C605 vdd.n42 iovss 0.91173f
C606 vdd.n52 iovss 0.6924f
C607 vdd.n54 iovss 0.60177f
C608 vdd.n55 iovss 0.55436f
C609 p2c.t0 iovss 0.2206f
C610 p2c.t1 iovss 0.45472f
C611 p2c.n1 iovss 0.21646f
C612 p2c.n2 iovss 0.75346f
C613 p2c.n3 iovss 1.9316f
.ends

