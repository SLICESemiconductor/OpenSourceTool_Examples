* NGSPICE file created from OTA_final.ext - technology: ihp-sg13g2

.subckt OTA_final ibias vinn vinp vout vdda vssa
X0 vssa vssa vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=44.7395p ps=0.39066m w=1u l=2u
X1 w_833_2071.t42 ibias.t12 vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X2 a_610_6649.t15 vinp.t0 w_833_2071.t45 w_833_2071.t19 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X3 w_833_2071.t21 vinn.t0 vout.t9 w_833_2071.t4 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X4 a_610_6649.t14 vinp.t1 w_833_2071.t18 w_833_2071.t30 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X5 vdda vdda vdda vdda sg13_lv_pmos ad=0.34p pd=2.68u as=81.07089p ps=0.63235m w=1u l=1u
X6 vdda a_610_6649.t28 vout.t3 vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X7 w_833_2071.t43 ibias.t13 vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X8 w_833_2071.t81 w_833_2071.t138 w_833_2071.t81 w_833_2071.t19 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X9 w_833_2071.t20 vinn.t1 vout.t16 w_833_2071.t56 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X10 vdda vdda vdda vdda sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X11 w_833_2071.t50 vinn.t2 vout.t14 w_833_2071.t52 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X12 w_833_2071.t31 vinn.t3 vout.t5 w_833_2071.t17 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X13 w_833_2071.t81 w_833_2071.t136 w_833_2071.t81 w_833_2071.t4 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X14 w_833_2071.t81 w_833_2071.t134 w_833_2071.t81 w_833_2071.t30 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X15 a_610_6649.t12 vinp.t2 w_833_2071.t11 w_833_2071.t0 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X16 vdda a_610_6649.t27 a_610_6649.t21 vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X17 w_833_2071.t75 w_833_2071.t132 w_833_2071.t75 w_833_2071.t56 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X18 vssa vssa vssa vssa sg13_lv_nmos ad=0.36p pd=2.72u as=0 ps=0 w=1u l=1u
X19 w_833_2071.t75 w_833_2071.t130 w_833_2071.t75 w_833_2071.t17 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X20 ibias.t10 ibias.t11 vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X21 w_833_2071.t75 w_833_2071.t128 w_833_2071.t75 w_833_2071.t0 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X22 vdda vdda vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X23 w_833_2071.t45 vinp.t3 a_610_6649.t8 w_833_2071.t56 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X24 vdda a_610_6649.t26 a_610_6649.t23 vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X25 w_833_2071.t18 vinp.t4 a_610_6649.t15 w_833_2071.t17 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X26 vdda vdda vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X27 a_610_6649.t13 vinp.t5 w_833_2071.t8 w_833_2071.t6 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X28 vout.t18 vinn.t4 w_833_2071.t21 w_833_2071.t0 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X29 w_833_2071.t44 vinp.t6 a_610_6649.t7 w_833_2071.t52 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X30 vdda a_610_6649.t29 vout.t2 vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X31 vssa vssa vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X32 vssa ibias.t14 w_833_2071.t43 vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X33 w_833_2071.t81 w_833_2071.t126 w_833_2071.t81 w_833_2071.t56 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X34 vssa vssa vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X35 vdda vdda vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X36 vdda a_610_6649.t30 vout.t1 vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X37 w_833_2071.t81 w_833_2071.t124 w_833_2071.t81 w_833_2071.t17 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X38 vssa vssa vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X39 vssa ibias.t9 ibias.t10 vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X40 w_833_2071.t81 w_833_2071.t122 w_833_2071.t81 w_833_2071.t0 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X41 vssa vssa vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X42 vdda a_610_6649.t25 a_610_6649.t17 vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X43 vdda vdda vdda vdda sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X44 vssa vssa vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X45 w_833_2071.t40 ibias.t15 vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X46 vdda vdda vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X47 vout.t17 vinn.t5 w_833_2071.t26 w_833_2071.t6 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X48 vdda a_610_6649.t24 a_610_6649.t19 vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X49 w_833_2071.t8 vinp.t7 a_610_6649.t6 w_833_2071.t24 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X50 vssa vssa vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X51 w_833_2071.t41 ibias.t16 vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X52 vdda vdda vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X53 vssa ibias.t17 w_833_2071.t42 vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X54 vdda a_610_6649.t31 vout.t0 vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X55 vssa vssa vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X56 w_833_2071.t10 vinn.t6 vout.t4 w_833_2071.t52 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X57 vssa vssa vssa vssa sg13_lv_nmos ad=0.36p pd=2.72u as=0 ps=0 w=1u l=1u
X58 vdda vdda vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X59 w_833_2071.t75 w_833_2071.t120 w_833_2071.t75 w_833_2071.t52 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X60 vout.t12 vinn.t7 w_833_2071.t60 w_833_2071.t15 sg13_lv_nmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.5u
X61 vssa vssa vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X62 w_833_2071.t26 vinn.t8 vout.t6 w_833_2071.t24 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X63 vdda vdda vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X64 w_833_2071.t33 vinn.t9 vout.t19 w_833_2071.t28 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X65 w_833_2071.t53 vinp.t8 a_610_6649.t14 w_833_2071.t52 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X66 a_610_6649.t11 vinp.t9 w_833_2071.t61 w_833_2071.t23 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X67 vssa ibias.t18 w_833_2071.t41 vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X68 a_610_6649.t5 vinp.t10 w_833_2071.t7 w_833_2071.t6 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X69 vssa vssa vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X70 w_833_2071.t81 w_833_2071.t118 w_833_2071.t81 w_833_2071.t52 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X71 vssa vssa vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X72 vdda vdda vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X73 ibias.t7 ibias.t8 vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X74 w_833_2071.t75 w_833_2071.t116 w_833_2071.t75 w_833_2071.t6 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X75 a_610_6649.t23 a_610_6649.t22 vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X76 a_610_6649.t2 vinp.t11 w_833_2071.t29 w_833_2071.t15 sg13_lv_nmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.5u
X77 vdda vdda vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X78 vssa vssa vssa vssa sg13_lv_nmos ad=0.36p pd=2.72u as=0 ps=0 w=1u l=1u
X79 vout.t8 vinn.t10 w_833_2071.t25 w_833_2071.t6 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X80 w_833_2071.t3 vinp.t12 a_610_6649.t10 w_833_2071.t28 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X81 vdda vdda vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X82 vout.t19 vinn.t11 w_833_2071.t50 w_833_2071.t9 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X83 vout.t15 vinn.t12 w_833_2071.t13 w_833_2071.t23 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X84 a_610_6649.t9 vinp.t13 w_833_2071.t33 w_833_2071.t2 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X85 w_833_2071.t61 vinp.t14 a_610_6649.t13 w_833_2071.t12 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X86 vssa ibias.t19 w_833_2071.t40 vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X87 w_833_2071.t81 w_833_2071.t114 w_833_2071.t81 w_833_2071.t6 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X88 w_833_2071.t7 vinp.t15 a_610_6649.t12 w_833_2071.t24 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X89 w_833_2071.t39 vinp.t16 a_610_6649.t11 w_833_2071.t38 sg13_lv_nmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.5u
X90 vssa ibias.t6 ibias.t7 vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X91 vssa vssa vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X92 vdda vdda vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X93 a_610_6649.t21 a_610_6649.t20 vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X94 w_833_2071.t75 w_833_2071.t112 w_833_2071.t75 w_833_2071.t24 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X95 vssa vssa vssa vssa sg13_lv_nmos ad=0.36p pd=2.72u as=0 ps=0 w=1u l=1u
X96 a_610_6649.t19 a_610_6649.t18 vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X97 vdda vdda vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X98 vout.t3 a_610_6649.t32 vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X99 w_833_2071.t25 vinn.t13 vout.t18 w_833_2071.t24 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X100 a_610_6649.t10 vinp.t17 w_833_2071.t44 w_833_2071.t9 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X101 vssa vssa vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X102 w_833_2071.t13 vinn.t14 vout.t17 w_833_2071.t12 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X103 vout.t13 vinn.t15 w_833_2071.t3 w_833_2071.t2 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X104 vdda vdda vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X105 vout.t11 vinn.t16 w_833_2071.t57 w_833_2071.t19 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X106 vout.t16 vinn.t17 w_833_2071.t27 w_833_2071.t15 sg13_lv_nmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.5u
X107 w_833_2071.t49 vinn.t18 vout.t15 w_833_2071.t38 sg13_lv_nmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.5u
X108 vout.t14 vinn.t19 w_833_2071.t32 w_833_2071.t30 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X109 w_833_2071.t1 vinp.t18 a_610_6649.t9 w_833_2071.t4 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X110 w_833_2071.t81 w_833_2071.t110 w_833_2071.t81 w_833_2071.t24 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X111 w_833_2071.t22 vinn.t20 vout.t10 w_833_2071.t28 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X112 vssa vssa vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X113 vssa vssa vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X114 a_610_6649.t4 vinp.t19 w_833_2071.t36 w_833_2071.t23 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X115 vdda vdda vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X116 w_833_2071.t109 w_833_2071.t107 w_833_2071.t75 w_833_2071.t15 sg13_lv_nmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=0.5u
X117 w_833_2071.t75 w_833_2071.t105 w_833_2071.t75 w_833_2071.t28 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X118 ibias.t4 ibias.t5 vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X119 a_610_6649.t17 a_610_6649.t16 vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X120 vssa vssa vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X121 w_833_2071.t75 w_833_2071.t103 w_833_2071.t75 w_833_2071.t23 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X122 vdda vdda vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X123 a_610_6649.t8 vinp.t20 w_833_2071.t16 w_833_2071.t15 sg13_lv_nmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.5u
X124 w_833_2071.t14 vinp.t21 a_610_6649.t3 w_833_2071.t28 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X125 vout.t2 a_610_6649.t33 vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X126 a_610_6649.t1 vinp.t22 w_833_2071.t63 w_833_2071.t19 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X127 a_610_6649.t7 vinp.t23 w_833_2071.t35 w_833_2071.t30 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X128 vssa vssa vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X129 vout.t7 vinn.t21 w_833_2071.t34 w_833_2071.t23 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X130 w_833_2071.t5 vinn.t22 vout.t13 w_833_2071.t4 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X131 w_833_2071.t57 vinn.t23 vout.t12 w_833_2071.t56 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X132 w_833_2071.t32 vinn.t24 vout.t11 w_833_2071.t17 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X133 w_833_2071.t102 w_833_2071.t100 w_833_2071.t81 w_833_2071.t15 sg13_lv_nmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=0.5u
X134 w_833_2071.t81 w_833_2071.t98 w_833_2071.t81 w_833_2071.t28 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X135 vout.t10 vinn.t25 w_833_2071.t10 w_833_2071.t9 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X136 vdda vdda vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X137 a_610_6649.t6 vinp.t24 w_833_2071.t1 w_833_2071.t0 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X138 w_833_2071.t36 vinp.t25 a_610_6649.t5 w_833_2071.t12 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X139 a_610_6649.t0 vinp.t26 w_833_2071.t22 w_833_2071.t2 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X140 vout.t1 a_610_6649.t34 vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X141 vssa ibias.t3 ibias.t4 vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X142 w_833_2071.t81 w_833_2071.t96 w_833_2071.t81 w_833_2071.t23 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X143 w_833_2071.t146 vinp.t27 a_610_6649.t4 w_833_2071.t38 sg13_lv_nmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.5u
X144 vdda vdda vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X145 w_833_2071.t75 w_833_2071.t94 w_833_2071.t75 w_833_2071.t9 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X146 w_833_2071.t75 w_833_2071.t92 w_833_2071.t75 w_833_2071.t2 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X147 w_833_2071.t75 w_833_2071.t90 w_833_2071.t75 w_833_2071.t12 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X148 ibias.t1 ibias.t2 vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X149 w_833_2071.t75 w_833_2071.t88 w_833_2071.t75 w_833_2071.t38 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X150 vssa vssa vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X151 a_610_6649.t3 vinp.t28 w_833_2071.t53 w_833_2071.t9 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X152 w_833_2071.t63 vinp.t29 a_610_6649.t2 w_833_2071.t56 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X153 vout.t9 vinn.t26 w_833_2071.t14 w_833_2071.t2 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X154 w_833_2071.t35 vinp.t30 a_610_6649.t1 w_833_2071.t17 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X155 w_833_2071.t34 vinn.t27 vout.t8 w_833_2071.t12 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X156 w_833_2071.t145 vinn.t28 vout.t7 w_833_2071.t38 sg13_lv_nmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.5u
X157 vdda vdda vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X158 vout.t6 vinn.t29 w_833_2071.t5 w_833_2071.t0 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X159 vdda vdda vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X160 vdda vdda vdda vdda sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X161 w_833_2071.t81 w_833_2071.t86 w_833_2071.t81 w_833_2071.t9 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X162 vout.t5 vinn.t30 w_833_2071.t20 w_833_2071.t19 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X163 vout.t4 vinn.t31 w_833_2071.t31 w_833_2071.t30 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X164 vssa vssa vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X165 w_833_2071.t81 w_833_2071.t84 w_833_2071.t81 w_833_2071.t12 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X166 w_833_2071.t81 w_833_2071.t82 w_833_2071.t81 w_833_2071.t2 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X167 w_833_2071.t11 vinp.t31 a_610_6649.t0 w_833_2071.t4 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X168 vssa ibias.t0 ibias.t1 vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X169 w_833_2071.t81 w_833_2071.t80 w_833_2071.t81 w_833_2071.t38 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X170 vout.t0 a_610_6649.t35 vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X171 vdda vdda vdda vdda sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X172 vssa vssa vssa vssa sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X173 w_833_2071.t75 w_833_2071.t78 w_833_2071.t75 w_833_2071.t19 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X174 w_833_2071.t75 w_833_2071.t76 w_833_2071.t75 w_833_2071.t30 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X175 w_833_2071.t75 w_833_2071.t74 w_833_2071.t75 w_833_2071.t4 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
R0 ibias.n22 ibias.n0 10.8172
R1 ibias.n22 ibias.n21 9.37277
R2 ibias.n15 ibias.t10 5.6534
R3 ibias.n20 ibias.t4 5.6534
R4 ibias.n10 ibias.t7 5.6534
R5 ibias.n5 ibias.t1 5.6534
R6 ibias.n11 ibias.t16 4.42794
R7 ibias.n13 ibias.t19 4.42666
R8 ibias.n3 ibias.t17 4.42666
R9 ibias.n1 ibias.t13 4.42557
R10 ibias ibias.n22 3.81636
R11 ibias.n21 ibias.n10 3.73245
R12 ibias.n5 ibias.n0 3.73245
R13 ibias.n15 ibias.n0 3.04514
R14 ibias.n21 ibias.n20 3.04514
R15 ibias.n2 ibias.t8 2.82253
R16 ibias.n1 ibias.t14 2.82253
R17 ibias.n13 ibias.t15 2.82253
R18 ibias.n14 ibias.t9 2.82253
R19 ibias.n12 ibias.t5 2.82253
R20 ibias.n11 ibias.t18 2.82253
R21 ibias.n17 ibias.t11 2.82253
R22 ibias.n18 ibias.t3 2.82253
R23 ibias.n7 ibias.t2 2.82253
R24 ibias.n8 ibias.t6 2.82253
R25 ibias.n3 ibias.t12 2.82253
R26 ibias.n4 ibias.t0 2.82253
R27 ibias.n2 ibias.n1 1.60563
R28 ibias.n14 ibias.n13 1.60563
R29 ibias.n12 ibias.n11 1.60563
R30 ibias.n18 ibias.n17 1.60563
R31 ibias.n8 ibias.n7 1.60563
R32 ibias.n4 ibias.n3 1.60563
R33 ibias.n16 ibias.n14 0.704016
R34 ibias.n19 ibias.n18 0.704016
R35 ibias.n9 ibias.n8 0.704016
R36 ibias.n6 ibias.n4 0.704016
R37 ibias.n9 ibias.n2 0.702736
R38 ibias.n19 ibias.n12 0.702736
R39 ibias.n17 ibias.n16 0.702736
R40 ibias.n7 ibias.n6 0.702736
R41 ibias.n16 ibias.n15 0.26531
R42 ibias.n20 ibias.n19 0.26531
R43 ibias.n10 ibias.n9 0.26531
R44 ibias.n6 ibias.n5 0.26531
R45 w_833_2071.n290 w_833_2071.n30 60.1886
R46 w_833_2071.n273 w_833_2071.t38 56.4268
R47 w_833_2071.n274 w_833_2071.n50 56.4268
R48 w_833_2071.n275 w_833_2071.n49 56.4268
R49 w_833_2071.n271 w_833_2071.n3 56.4268
R50 w_833_2071.n270 w_833_2071.n6 56.4268
R51 w_833_2071.n269 w_833_2071.n7 56.4268
R52 w_833_2071.n278 w_833_2071.n46 56.4268
R53 w_833_2071.n279 w_833_2071.n45 56.4268
R54 w_833_2071.n267 w_833_2071.n9 56.4268
R55 w_833_2071.n280 w_833_2071.n44 56.4268
R56 w_833_2071.n266 w_833_2071.n10 56.4268
R57 w_833_2071.n265 w_833_2071.n11 56.4268
R58 w_833_2071.n282 w_833_2071.n42 56.4268
R59 w_833_2071.n283 w_833_2071.n41 56.4268
R60 w_833_2071.n284 w_833_2071.n40 56.4268
R61 w_833_2071.n261 w_833_2071.n15 56.4268
R62 w_833_2071.n260 w_833_2071.n16 56.4268
R63 w_833_2071.t52 w_833_2071.n38 56.4268
R64 w_833_2071.n259 w_833_2071.n17 56.4268
R65 w_833_2071.n286 w_833_2071.n34 56.4268
R66 w_833_2071.n287 w_833_2071.n33 56.4268
R67 w_833_2071.n257 w_833_2071.n19 56.4268
R68 w_833_2071.n256 w_833_2071.n21 56.4268
R69 w_833_2071.n255 w_833_2071.n22 56.4268
R70 w_833_2071.n291 w_833_2071.n27 56.4268
R71 w_833_2071.n292 w_833_2071.n26 56.4268
R72 w_833_2071.n288 w_833_2071.t17 52.6651
R73 w_833_2071.t6 w_833_2071.n47 48.9033
R74 w_833_2071.n263 w_833_2071.t2 48.9033
R75 w_833_2071.t15 w_833_2071.n24 48.9033
R76 w_833_2071.n276 w_833_2071.t12 45.1416
R77 w_833_2071.t28 w_833_2071.n13 45.1416
R78 w_833_2071.n254 w_833_2071.t56 45.1416
R79 w_833_2071.t19 w_833_2071.n31 41.3798
R80 w_833_2071.t23 w_833_2071.n2 37.6181
R81 w_833_2071.n285 w_833_2071.t9 37.6181
R82 w_833_2071.n268 w_833_2071.t24 33.8563
R83 w_833_2071.t4 w_833_2071.n43 33.8563
R84 w_833_2071.t30 w_833_2071.n18 30.0945
R85 w_833_2071.n258 w_833_2071.t30 26.3328
R86 w_833_2071.t24 w_833_2071.n8 22.571
R87 w_833_2071.n281 w_833_2071.t4 22.571
R88 w_833_2071.n272 w_833_2071.t23 18.8093
R89 w_833_2071.t9 w_833_2071.n39 18.8093
R90 w_833_2071.n53 w_833_2071.t38 17.3178
R91 w_833_2071.t75 w_833_2071.n94 17.0005
R92 w_833_2071.n56 w_833_2071.n25 17.0005
R93 w_833_2071.n56 w_833_2071.n26 17.0005
R94 w_833_2071.n56 w_833_2071.n24 17.0005
R95 w_833_2071.n56 w_833_2071.n27 17.0005
R96 w_833_2071.n56 w_833_2071.n23 17.0005
R97 w_833_2071.n56 w_833_2071.n30 17.0005
R98 w_833_2071.n56 w_833_2071.n22 17.0005
R99 w_833_2071.n56 w_833_2071.n31 17.0005
R100 w_833_2071.n56 w_833_2071.n21 17.0005
R101 w_833_2071.n56 w_833_2071.n32 17.0005
R102 w_833_2071.n56 w_833_2071.n19 17.0005
R103 w_833_2071.n56 w_833_2071.n33 17.0005
R104 w_833_2071.n56 w_833_2071.n18 17.0005
R105 w_833_2071.n56 w_833_2071.n34 17.0005
R106 w_833_2071.n56 w_833_2071.n17 17.0005
R107 w_833_2071.n56 w_833_2071.n38 17.0005
R108 w_833_2071.n56 w_833_2071.n16 17.0005
R109 w_833_2071.n56 w_833_2071.n39 17.0005
R110 w_833_2071.n56 w_833_2071.n15 17.0005
R111 w_833_2071.n56 w_833_2071.n40 17.0005
R112 w_833_2071.n56 w_833_2071.n13 17.0005
R113 w_833_2071.n56 w_833_2071.n41 17.0005
R114 w_833_2071.n56 w_833_2071.n12 17.0005
R115 w_833_2071.n56 w_833_2071.n42 17.0005
R116 w_833_2071.n56 w_833_2071.n11 17.0005
R117 w_833_2071.n56 w_833_2071.n43 17.0005
R118 w_833_2071.n56 w_833_2071.n10 17.0005
R119 w_833_2071.n56 w_833_2071.n44 17.0005
R120 w_833_2071.n56 w_833_2071.n9 17.0005
R121 w_833_2071.n56 w_833_2071.n45 17.0005
R122 w_833_2071.n56 w_833_2071.n8 17.0005
R123 w_833_2071.n56 w_833_2071.n46 17.0005
R124 w_833_2071.n56 w_833_2071.n7 17.0005
R125 w_833_2071.n56 w_833_2071.n47 17.0005
R126 w_833_2071.n56 w_833_2071.n6 17.0005
R127 w_833_2071.n56 w_833_2071.n48 17.0005
R128 w_833_2071.n56 w_833_2071.n3 17.0005
R129 w_833_2071.n56 w_833_2071.n49 17.0005
R130 w_833_2071.n56 w_833_2071.n2 17.0005
R131 w_833_2071.n56 w_833_2071.n50 17.0005
R132 w_833_2071.n56 w_833_2071.t38 17.0005
R133 w_833_2071.n326 w_833_2071.n56 17.0005
R134 w_833_2071.n54 w_833_2071.n25 17.0005
R135 w_833_2071.n54 w_833_2071.n26 17.0005
R136 w_833_2071.n54 w_833_2071.n24 17.0005
R137 w_833_2071.n54 w_833_2071.n27 17.0005
R138 w_833_2071.n54 w_833_2071.n23 17.0005
R139 w_833_2071.n54 w_833_2071.n30 17.0005
R140 w_833_2071.n54 w_833_2071.n22 17.0005
R141 w_833_2071.n54 w_833_2071.n31 17.0005
R142 w_833_2071.n54 w_833_2071.n21 17.0005
R143 w_833_2071.n54 w_833_2071.n32 17.0005
R144 w_833_2071.n54 w_833_2071.n19 17.0005
R145 w_833_2071.n54 w_833_2071.n33 17.0005
R146 w_833_2071.n54 w_833_2071.n18 17.0005
R147 w_833_2071.n54 w_833_2071.n34 17.0005
R148 w_833_2071.n54 w_833_2071.n17 17.0005
R149 w_833_2071.n54 w_833_2071.n38 17.0005
R150 w_833_2071.n54 w_833_2071.n16 17.0005
R151 w_833_2071.n54 w_833_2071.n39 17.0005
R152 w_833_2071.n54 w_833_2071.n15 17.0005
R153 w_833_2071.n54 w_833_2071.n40 17.0005
R154 w_833_2071.n54 w_833_2071.n13 17.0005
R155 w_833_2071.n54 w_833_2071.n41 17.0005
R156 w_833_2071.n54 w_833_2071.n12 17.0005
R157 w_833_2071.n54 w_833_2071.n42 17.0005
R158 w_833_2071.n54 w_833_2071.n11 17.0005
R159 w_833_2071.n54 w_833_2071.n43 17.0005
R160 w_833_2071.n54 w_833_2071.n10 17.0005
R161 w_833_2071.n54 w_833_2071.n44 17.0005
R162 w_833_2071.n54 w_833_2071.n9 17.0005
R163 w_833_2071.n54 w_833_2071.n45 17.0005
R164 w_833_2071.n54 w_833_2071.n8 17.0005
R165 w_833_2071.n54 w_833_2071.n46 17.0005
R166 w_833_2071.n54 w_833_2071.n7 17.0005
R167 w_833_2071.n54 w_833_2071.n47 17.0005
R168 w_833_2071.n54 w_833_2071.n6 17.0005
R169 w_833_2071.n54 w_833_2071.n48 17.0005
R170 w_833_2071.n54 w_833_2071.n3 17.0005
R171 w_833_2071.n54 w_833_2071.n49 17.0005
R172 w_833_2071.n54 w_833_2071.n2 17.0005
R173 w_833_2071.n54 w_833_2071.n50 17.0005
R174 w_833_2071.n54 w_833_2071.t38 17.0005
R175 w_833_2071.n326 w_833_2071.n54 17.0005
R176 w_833_2071.n57 w_833_2071.n25 17.0005
R177 w_833_2071.n57 w_833_2071.n26 17.0005
R178 w_833_2071.n57 w_833_2071.n24 17.0005
R179 w_833_2071.n57 w_833_2071.n27 17.0005
R180 w_833_2071.n57 w_833_2071.n23 17.0005
R181 w_833_2071.n57 w_833_2071.n30 17.0005
R182 w_833_2071.n57 w_833_2071.n22 17.0005
R183 w_833_2071.n57 w_833_2071.n31 17.0005
R184 w_833_2071.n57 w_833_2071.n21 17.0005
R185 w_833_2071.n57 w_833_2071.n32 17.0005
R186 w_833_2071.n57 w_833_2071.n19 17.0005
R187 w_833_2071.n57 w_833_2071.n33 17.0005
R188 w_833_2071.n57 w_833_2071.n18 17.0005
R189 w_833_2071.n57 w_833_2071.n34 17.0005
R190 w_833_2071.n57 w_833_2071.n17 17.0005
R191 w_833_2071.n57 w_833_2071.n38 17.0005
R192 w_833_2071.n57 w_833_2071.n16 17.0005
R193 w_833_2071.n57 w_833_2071.n39 17.0005
R194 w_833_2071.n57 w_833_2071.n15 17.0005
R195 w_833_2071.n57 w_833_2071.n40 17.0005
R196 w_833_2071.n57 w_833_2071.n13 17.0005
R197 w_833_2071.n57 w_833_2071.n41 17.0005
R198 w_833_2071.n57 w_833_2071.n12 17.0005
R199 w_833_2071.n57 w_833_2071.n42 17.0005
R200 w_833_2071.n57 w_833_2071.n11 17.0005
R201 w_833_2071.n57 w_833_2071.n43 17.0005
R202 w_833_2071.n57 w_833_2071.n10 17.0005
R203 w_833_2071.n57 w_833_2071.n44 17.0005
R204 w_833_2071.n57 w_833_2071.n9 17.0005
R205 w_833_2071.n57 w_833_2071.n45 17.0005
R206 w_833_2071.n57 w_833_2071.n8 17.0005
R207 w_833_2071.n57 w_833_2071.n46 17.0005
R208 w_833_2071.n57 w_833_2071.n7 17.0005
R209 w_833_2071.n57 w_833_2071.n47 17.0005
R210 w_833_2071.n57 w_833_2071.n6 17.0005
R211 w_833_2071.n57 w_833_2071.n48 17.0005
R212 w_833_2071.n57 w_833_2071.n3 17.0005
R213 w_833_2071.n57 w_833_2071.n49 17.0005
R214 w_833_2071.n57 w_833_2071.n2 17.0005
R215 w_833_2071.n57 w_833_2071.n50 17.0005
R216 w_833_2071.n57 w_833_2071.t38 17.0005
R217 w_833_2071.n326 w_833_2071.n57 17.0005
R218 w_833_2071.n325 w_833_2071.n25 17.0005
R219 w_833_2071.n325 w_833_2071.n26 17.0005
R220 w_833_2071.n325 w_833_2071.n24 17.0005
R221 w_833_2071.n325 w_833_2071.n27 17.0005
R222 w_833_2071.n325 w_833_2071.n23 17.0005
R223 w_833_2071.n325 w_833_2071.n30 17.0005
R224 w_833_2071.n325 w_833_2071.n22 17.0005
R225 w_833_2071.n325 w_833_2071.n31 17.0005
R226 w_833_2071.n325 w_833_2071.n21 17.0005
R227 w_833_2071.n325 w_833_2071.n32 17.0005
R228 w_833_2071.n325 w_833_2071.n19 17.0005
R229 w_833_2071.n325 w_833_2071.n33 17.0005
R230 w_833_2071.n325 w_833_2071.n18 17.0005
R231 w_833_2071.n325 w_833_2071.n34 17.0005
R232 w_833_2071.n325 w_833_2071.n17 17.0005
R233 w_833_2071.n325 w_833_2071.n38 17.0005
R234 w_833_2071.n325 w_833_2071.n16 17.0005
R235 w_833_2071.n325 w_833_2071.n39 17.0005
R236 w_833_2071.n325 w_833_2071.n15 17.0005
R237 w_833_2071.n325 w_833_2071.n40 17.0005
R238 w_833_2071.n325 w_833_2071.n13 17.0005
R239 w_833_2071.n325 w_833_2071.n41 17.0005
R240 w_833_2071.n325 w_833_2071.n12 17.0005
R241 w_833_2071.n325 w_833_2071.n42 17.0005
R242 w_833_2071.n325 w_833_2071.n11 17.0005
R243 w_833_2071.n325 w_833_2071.n43 17.0005
R244 w_833_2071.n325 w_833_2071.n10 17.0005
R245 w_833_2071.n325 w_833_2071.n44 17.0005
R246 w_833_2071.n325 w_833_2071.n9 17.0005
R247 w_833_2071.n325 w_833_2071.n45 17.0005
R248 w_833_2071.n325 w_833_2071.n8 17.0005
R249 w_833_2071.n325 w_833_2071.n46 17.0005
R250 w_833_2071.n325 w_833_2071.n7 17.0005
R251 w_833_2071.n325 w_833_2071.n47 17.0005
R252 w_833_2071.n325 w_833_2071.n6 17.0005
R253 w_833_2071.n325 w_833_2071.n48 17.0005
R254 w_833_2071.n325 w_833_2071.n3 17.0005
R255 w_833_2071.n325 w_833_2071.n49 17.0005
R256 w_833_2071.n325 w_833_2071.n2 17.0005
R257 w_833_2071.n325 w_833_2071.n50 17.0005
R258 w_833_2071.n325 w_833_2071.t38 17.0005
R259 w_833_2071.n326 w_833_2071.n325 17.0005
R260 w_833_2071.n293 w_833_2071.n273 17.0005
R261 w_833_2071.n293 w_833_2071.n274 17.0005
R262 w_833_2071.n293 w_833_2071.n272 17.0005
R263 w_833_2071.n293 w_833_2071.n275 17.0005
R264 w_833_2071.n293 w_833_2071.n271 17.0005
R265 w_833_2071.n293 w_833_2071.n276 17.0005
R266 w_833_2071.n293 w_833_2071.n270 17.0005
R267 w_833_2071.n293 w_833_2071.n277 17.0005
R268 w_833_2071.n293 w_833_2071.n269 17.0005
R269 w_833_2071.n293 w_833_2071.n278 17.0005
R270 w_833_2071.n293 w_833_2071.n268 17.0005
R271 w_833_2071.n293 w_833_2071.n279 17.0005
R272 w_833_2071.n293 w_833_2071.n267 17.0005
R273 w_833_2071.n293 w_833_2071.n280 17.0005
R274 w_833_2071.n293 w_833_2071.n266 17.0005
R275 w_833_2071.n293 w_833_2071.n281 17.0005
R276 w_833_2071.n293 w_833_2071.n265 17.0005
R277 w_833_2071.n293 w_833_2071.n282 17.0005
R278 w_833_2071.n293 w_833_2071.n263 17.0005
R279 w_833_2071.n293 w_833_2071.n283 17.0005
R280 w_833_2071.n293 w_833_2071.n262 17.0005
R281 w_833_2071.n293 w_833_2071.n284 17.0005
R282 w_833_2071.n293 w_833_2071.n261 17.0005
R283 w_833_2071.n293 w_833_2071.n285 17.0005
R284 w_833_2071.n293 w_833_2071.n260 17.0005
R285 w_833_2071.n293 w_833_2071.t52 17.0005
R286 w_833_2071.n293 w_833_2071.n259 17.0005
R287 w_833_2071.n293 w_833_2071.n286 17.0005
R288 w_833_2071.n293 w_833_2071.n258 17.0005
R289 w_833_2071.n293 w_833_2071.n287 17.0005
R290 w_833_2071.n293 w_833_2071.n257 17.0005
R291 w_833_2071.n293 w_833_2071.n288 17.0005
R292 w_833_2071.n293 w_833_2071.n256 17.0005
R293 w_833_2071.n293 w_833_2071.n289 17.0005
R294 w_833_2071.n293 w_833_2071.n255 17.0005
R295 w_833_2071.n293 w_833_2071.n290 17.0005
R296 w_833_2071.n293 w_833_2071.n254 17.0005
R297 w_833_2071.n293 w_833_2071.n291 17.0005
R298 w_833_2071.n293 w_833_2071.n253 17.0005
R299 w_833_2071.n293 w_833_2071.n292 17.0005
R300 w_833_2071.n194 w_833_2071.t81 17.0005
R301 w_833_2071.n55 w_833_2071.n26 17.0005
R302 w_833_2071.n55 w_833_2071.n24 17.0005
R303 w_833_2071.n55 w_833_2071.n27 17.0005
R304 w_833_2071.n55 w_833_2071.n23 17.0005
R305 w_833_2071.n55 w_833_2071.n30 17.0005
R306 w_833_2071.n55 w_833_2071.n22 17.0005
R307 w_833_2071.n55 w_833_2071.n31 17.0005
R308 w_833_2071.n55 w_833_2071.n21 17.0005
R309 w_833_2071.n55 w_833_2071.n32 17.0005
R310 w_833_2071.n55 w_833_2071.n19 17.0005
R311 w_833_2071.n55 w_833_2071.n33 17.0005
R312 w_833_2071.n55 w_833_2071.n18 17.0005
R313 w_833_2071.n55 w_833_2071.n34 17.0005
R314 w_833_2071.n55 w_833_2071.n17 17.0005
R315 w_833_2071.n55 w_833_2071.n38 17.0005
R316 w_833_2071.n55 w_833_2071.n16 17.0005
R317 w_833_2071.n55 w_833_2071.n39 17.0005
R318 w_833_2071.n55 w_833_2071.n15 17.0005
R319 w_833_2071.n142 w_833_2071.n55 17.0005
R320 w_833_2071.n55 w_833_2071.n25 17.0005
R321 w_833_2071.n326 w_833_2071.n55 17.0005
R322 w_833_2071.n55 w_833_2071.t38 17.0005
R323 w_833_2071.n55 w_833_2071.n50 17.0005
R324 w_833_2071.n55 w_833_2071.n2 17.0005
R325 w_833_2071.n55 w_833_2071.n49 17.0005
R326 w_833_2071.n55 w_833_2071.n3 17.0005
R327 w_833_2071.n55 w_833_2071.n48 17.0005
R328 w_833_2071.n55 w_833_2071.n6 17.0005
R329 w_833_2071.n55 w_833_2071.n47 17.0005
R330 w_833_2071.n55 w_833_2071.n7 17.0005
R331 w_833_2071.n55 w_833_2071.n46 17.0005
R332 w_833_2071.n55 w_833_2071.n8 17.0005
R333 w_833_2071.n55 w_833_2071.n45 17.0005
R334 w_833_2071.n55 w_833_2071.n9 17.0005
R335 w_833_2071.n55 w_833_2071.n44 17.0005
R336 w_833_2071.n55 w_833_2071.n10 17.0005
R337 w_833_2071.n55 w_833_2071.n43 17.0005
R338 w_833_2071.n55 w_833_2071.n11 17.0005
R339 w_833_2071.n55 w_833_2071.n42 17.0005
R340 w_833_2071.n55 w_833_2071.n12 17.0005
R341 w_833_2071.n55 w_833_2071.n41 17.0005
R342 w_833_2071.n55 w_833_2071.n13 17.0005
R343 w_833_2071.n55 w_833_2071.n40 17.0005
R344 w_833_2071.n327 w_833_2071.n25 17.0005
R345 w_833_2071.n327 w_833_2071.n26 17.0005
R346 w_833_2071.n327 w_833_2071.n24 17.0005
R347 w_833_2071.n327 w_833_2071.n27 17.0005
R348 w_833_2071.n327 w_833_2071.n23 17.0005
R349 w_833_2071.n327 w_833_2071.n30 17.0005
R350 w_833_2071.n327 w_833_2071.n22 17.0005
R351 w_833_2071.n327 w_833_2071.n31 17.0005
R352 w_833_2071.n327 w_833_2071.n21 17.0005
R353 w_833_2071.n327 w_833_2071.n32 17.0005
R354 w_833_2071.n327 w_833_2071.n19 17.0005
R355 w_833_2071.n327 w_833_2071.n33 17.0005
R356 w_833_2071.n327 w_833_2071.n18 17.0005
R357 w_833_2071.n327 w_833_2071.n34 17.0005
R358 w_833_2071.n327 w_833_2071.n17 17.0005
R359 w_833_2071.n327 w_833_2071.n38 17.0005
R360 w_833_2071.n327 w_833_2071.n16 17.0005
R361 w_833_2071.n327 w_833_2071.n39 17.0005
R362 w_833_2071.n327 w_833_2071.n15 17.0005
R363 w_833_2071.n327 w_833_2071.n40 17.0005
R364 w_833_2071.n327 w_833_2071.n13 17.0005
R365 w_833_2071.n327 w_833_2071.n41 17.0005
R366 w_833_2071.n327 w_833_2071.n12 17.0005
R367 w_833_2071.n327 w_833_2071.n42 17.0005
R368 w_833_2071.n327 w_833_2071.n11 17.0005
R369 w_833_2071.n327 w_833_2071.n43 17.0005
R370 w_833_2071.n327 w_833_2071.n10 17.0005
R371 w_833_2071.n327 w_833_2071.n44 17.0005
R372 w_833_2071.n327 w_833_2071.n9 17.0005
R373 w_833_2071.n327 w_833_2071.n45 17.0005
R374 w_833_2071.n327 w_833_2071.n8 17.0005
R375 w_833_2071.n327 w_833_2071.n46 17.0005
R376 w_833_2071.n327 w_833_2071.n7 17.0005
R377 w_833_2071.n327 w_833_2071.n47 17.0005
R378 w_833_2071.n327 w_833_2071.n6 17.0005
R379 w_833_2071.n327 w_833_2071.n48 17.0005
R380 w_833_2071.n327 w_833_2071.n3 17.0005
R381 w_833_2071.n327 w_833_2071.n49 17.0005
R382 w_833_2071.n327 w_833_2071.n2 17.0005
R383 w_833_2071.n327 w_833_2071.n50 17.0005
R384 w_833_2071.n327 w_833_2071.t38 17.0005
R385 w_833_2071.n327 w_833_2071.n326 17.0005
R386 w_833_2071.n175 w_833_2071.t42 15.3683
R387 w_833_2071.n139 w_833_2071.t43 15.3683
R388 w_833_2071.n289 w_833_2071.t19 15.0475
R389 w_833_2071.n104 w_833_2071.t103 15.0005
R390 w_833_2071.n106 w_833_2071.t90 15.0005
R391 w_833_2071.n107 w_833_2071.t116 15.0005
R392 w_833_2071.n319 w_833_2071.t112 15.0005
R393 w_833_2071.n317 w_833_2071.t128 15.0005
R394 w_833_2071.n315 w_833_2071.t74 15.0005
R395 w_833_2071.n313 w_833_2071.t92 15.0005
R396 w_833_2071.n311 w_833_2071.t105 15.0005
R397 w_833_2071.n309 w_833_2071.t94 15.0005
R398 w_833_2071.n307 w_833_2071.t120 15.0005
R399 w_833_2071.n305 w_833_2071.t76 15.0005
R400 w_833_2071.n303 w_833_2071.t130 15.0005
R401 w_833_2071.n301 w_833_2071.t78 15.0005
R402 w_833_2071.n299 w_833_2071.t132 15.0005
R403 w_833_2071.n297 w_833_2071.t107 15.0005
R404 w_833_2071.n102 w_833_2071.t88 15.0005
R405 w_833_2071.n173 w_833_2071.t80 15.0005
R406 w_833_2071.n171 w_833_2071.t96 15.0005
R407 w_833_2071.n169 w_833_2071.t84 15.0005
R408 w_833_2071.n168 w_833_2071.t114 15.0005
R409 w_833_2071.n166 w_833_2071.t110 15.0005
R410 w_833_2071.n164 w_833_2071.t122 15.0005
R411 w_833_2071.n162 w_833_2071.t136 15.0005
R412 w_833_2071.n160 w_833_2071.t82 15.0005
R413 w_833_2071.n158 w_833_2071.t98 15.0005
R414 w_833_2071.n156 w_833_2071.t86 15.0005
R415 w_833_2071.n154 w_833_2071.t118 15.0005
R416 w_833_2071.n152 w_833_2071.t134 15.0005
R417 w_833_2071.n150 w_833_2071.t124 15.0005
R418 w_833_2071.n148 w_833_2071.t138 15.0005
R419 w_833_2071.n146 w_833_2071.t126 15.0005
R420 w_833_2071.n144 w_833_2071.t100 15.0005
R421 w_833_2071.n175 w_833_2071.t40 14.6976
R422 w_833_2071.n139 w_833_2071.t41 14.6976
R423 w_833_2071.n326 w_833_2071.n53 14.1283
R424 w_833_2071.n252 w_833_2071.n251 13.8647
R425 w_833_2071.n247 w_833_2071.n246 13.5377
R426 w_833_2071.n230 w_833_2071.n229 13.5377
R427 w_833_2071.n213 w_833_2071.n212 13.5377
R428 w_833_2071.n249 w_833_2071.n248 13.5377
R429 w_833_2071.n196 w_833_2071.n195 13.5005
R430 w_833_2071.n251 w_833_2071.n250 13.5005
R431 w_833_2071.t12 w_833_2071.n48 11.2858
R432 w_833_2071.n262 w_833_2071.t28 11.2858
R433 w_833_2071.t56 w_833_2071.n23 11.2858
R434 w_833_2071.n141 w_833_2071.n140 9.0005
R435 w_833_2071.n183 w_833_2071.n108 9.0005
R436 w_833_2071.n177 w_833_2071.n176 9.0005
R437 w_833_2071.n325 w_833_2071.n68 8.46995
R438 w_833_2071.n325 w_833_2071.n64 8.46995
R439 w_833_2071.n325 w_833_2071.n62 8.46995
R440 w_833_2071.n325 w_833_2071.n71 8.46995
R441 w_833_2071.n325 w_833_2071.n60 8.46995
R442 w_833_2071.n325 w_833_2071.n58 8.46995
R443 w_833_2071.n138 w_833_2071.n55 8.46995
R444 w_833_2071.n130 w_833_2071.n55 8.46995
R445 w_833_2071.n180 w_833_2071.n55 8.46995
R446 w_833_2071.n190 w_833_2071.n55 8.46995
R447 w_833_2071.n186 w_833_2071.n55 8.46995
R448 w_833_2071.n124 w_833_2071.n55 8.46995
R449 w_833_2071.n134 w_833_2071.n55 8.46995
R450 w_833_2071.t75 w_833_2071.n92 8.46336
R451 w_833_2071.t81 w_833_2071.n109 8.45649
R452 w_833_2071.n273 w_833_2071.n50 7.52401
R453 w_833_2071.n274 w_833_2071.n2 7.52401
R454 w_833_2071.n272 w_833_2071.n49 7.52401
R455 w_833_2071.n275 w_833_2071.n3 7.52401
R456 w_833_2071.n271 w_833_2071.n48 7.52401
R457 w_833_2071.n276 w_833_2071.n6 7.52401
R458 w_833_2071.n270 w_833_2071.n47 7.52401
R459 w_833_2071.n277 w_833_2071.t6 7.52401
R460 w_833_2071.n277 w_833_2071.n7 7.52401
R461 w_833_2071.n269 w_833_2071.n46 7.52401
R462 w_833_2071.n278 w_833_2071.n8 7.52401
R463 w_833_2071.n268 w_833_2071.n45 7.52401
R464 w_833_2071.n279 w_833_2071.n9 7.52401
R465 w_833_2071.n280 w_833_2071.n10 7.52401
R466 w_833_2071.n266 w_833_2071.n43 7.52401
R467 w_833_2071.n281 w_833_2071.n11 7.52401
R468 w_833_2071.n265 w_833_2071.n42 7.52401
R469 w_833_2071.n282 w_833_2071.n12 7.52401
R470 w_833_2071.t2 w_833_2071.n12 7.52401
R471 w_833_2071.n263 w_833_2071.n41 7.52401
R472 w_833_2071.n283 w_833_2071.n13 7.52401
R473 w_833_2071.n262 w_833_2071.n40 7.52401
R474 w_833_2071.n284 w_833_2071.n15 7.52401
R475 w_833_2071.n261 w_833_2071.n39 7.52401
R476 w_833_2071.n285 w_833_2071.n16 7.52401
R477 w_833_2071.n260 w_833_2071.n38 7.52401
R478 w_833_2071.t52 w_833_2071.n17 7.52401
R479 w_833_2071.n259 w_833_2071.n34 7.52401
R480 w_833_2071.n286 w_833_2071.n18 7.52401
R481 w_833_2071.n258 w_833_2071.n33 7.52401
R482 w_833_2071.n287 w_833_2071.n19 7.52401
R483 w_833_2071.n257 w_833_2071.n32 7.52401
R484 w_833_2071.n288 w_833_2071.n21 7.52401
R485 w_833_2071.n256 w_833_2071.n31 7.52401
R486 w_833_2071.n289 w_833_2071.n22 7.52401
R487 w_833_2071.n255 w_833_2071.n30 7.52401
R488 w_833_2071.n290 w_833_2071.n23 7.52401
R489 w_833_2071.n254 w_833_2071.n27 7.52401
R490 w_833_2071.n291 w_833_2071.n24 7.52401
R491 w_833_2071.n253 w_833_2071.t15 7.52401
R492 w_833_2071.n253 w_833_2071.n26 7.52401
R493 w_833_2071.n292 w_833_2071.n25 7.52401
R494 w_833_2071.n238 w_833_2071.t29 6.43891
R495 w_833_2071.n221 w_833_2071.t27 6.43891
R496 w_833_2071.n204 w_833_2071.t16 6.43891
R497 w_833_2071.n29 w_833_2071.t60 6.43891
R498 w_833_2071.n52 w_833_2071.t39 6.4061
R499 w_833_2071.n231 w_833_2071.t49 6.4061
R500 w_833_2071.n214 w_833_2071.t146 6.4061
R501 w_833_2071.n197 w_833_2071.t145 6.4061
R502 w_833_2071.n176 w_833_2071.n175 6.15663
R503 w_833_2071.n140 w_833_2071.n139 6.15663
R504 w_833_2071.n51 w_833_2071.t61 6.12323
R505 w_833_2071.n4 w_833_2071.t8 6.12323
R506 w_833_2071.n232 w_833_2071.t13 6.12323
R507 w_833_2071.n234 w_833_2071.t26 6.12323
R508 w_833_2071.n236 w_833_2071.t5 6.12323
R509 w_833_2071.n243 w_833_2071.t44 6.12323
R510 w_833_2071.n241 w_833_2071.t35 6.12323
R511 w_833_2071.n239 w_833_2071.t63 6.12323
R512 w_833_2071.n215 w_833_2071.t36 6.12323
R513 w_833_2071.n217 w_833_2071.t7 6.12323
R514 w_833_2071.n219 w_833_2071.t11 6.12323
R515 w_833_2071.n226 w_833_2071.t10 6.12323
R516 w_833_2071.n224 w_833_2071.t31 6.12323
R517 w_833_2071.n222 w_833_2071.t20 6.12323
R518 w_833_2071.n198 w_833_2071.t34 6.12323
R519 w_833_2071.n200 w_833_2071.t25 6.12323
R520 w_833_2071.n202 w_833_2071.t21 6.12323
R521 w_833_2071.n209 w_833_2071.t53 6.12323
R522 w_833_2071.n207 w_833_2071.t18 6.12323
R523 w_833_2071.n205 w_833_2071.t45 6.12323
R524 w_833_2071.n36 w_833_2071.t50 6.12323
R525 w_833_2071.n35 w_833_2071.t32 6.12323
R526 w_833_2071.n28 w_833_2071.t57 6.12323
R527 w_833_2071.t75 w_833_2071.n322 6.12223
R528 w_833_2071.t81 w_833_2071.n193 6.12223
R529 w_833_2071.t1 w_833_2071.n329 6.12223
R530 w_833_2071.n246 w_833_2071.t3 5.67005
R531 w_833_2071.n229 w_833_2071.t22 5.67005
R532 w_833_2071.n212 w_833_2071.t14 5.67005
R533 w_833_2071.n248 w_833_2071.t33 5.67005
R534 w_833_2071.n325 w_833_2071.n66 5.61281
R535 w_833_2071.n325 w_833_2071.n65 5.61281
R536 w_833_2071.n325 w_833_2071.n69 5.61281
R537 w_833_2071.n325 w_833_2071.n63 5.61281
R538 w_833_2071.n325 w_833_2071.n70 5.61281
R539 w_833_2071.n325 w_833_2071.n61 5.61281
R540 w_833_2071.n325 w_833_2071.n72 5.61281
R541 w_833_2071.n325 w_833_2071.n59 5.61281
R542 w_833_2071.n325 w_833_2071.n324 5.61281
R543 w_833_2071.n178 w_833_2071.n55 5.61281
R544 w_833_2071.n182 w_833_2071.n55 5.61281
R545 w_833_2071.n192 w_833_2071.n55 5.61281
R546 w_833_2071.n188 w_833_2071.n55 5.61281
R547 w_833_2071.n184 w_833_2071.n55 5.61281
R548 w_833_2071.n132 w_833_2071.n55 5.61281
R549 w_833_2071.n128 w_833_2071.n55 5.61281
R550 w_833_2071.n126 w_833_2071.n55 5.61281
R551 w_833_2071.n325 w_833_2071.n67 5.61121
R552 w_833_2071.n136 w_833_2071.n55 5.61121
R553 w_833_2071.n323 w_833_2071.t75 5.56245
R554 w_833_2071.t75 w_833_2071.n79 5.56245
R555 w_833_2071.t75 w_833_2071.n81 5.56245
R556 w_833_2071.t75 w_833_2071.n83 5.56245
R557 w_833_2071.t75 w_833_2071.n85 5.56245
R558 w_833_2071.t75 w_833_2071.n87 5.56245
R559 w_833_2071.t75 w_833_2071.n89 5.56245
R560 w_833_2071.t75 w_833_2071.n91 5.56245
R561 w_833_2071.t75 w_833_2071.n96 5.56245
R562 w_833_2071.t75 w_833_2071.n98 5.56245
R563 w_833_2071.t75 w_833_2071.n100 5.56245
R564 w_833_2071.t75 w_833_2071.n321 5.56245
R565 w_833_2071.t75 w_833_2071.n77 5.56245
R566 w_833_2071.t75 w_833_2071.n75 5.56245
R567 w_833_2071.n295 w_833_2071.t109 5.56245
R568 w_833_2071.t81 w_833_2071.n121 5.56245
R569 w_833_2071.t81 w_833_2071.n120 5.56245
R570 w_833_2071.t81 w_833_2071.n119 5.56245
R571 w_833_2071.t81 w_833_2071.n118 5.56245
R572 w_833_2071.t81 w_833_2071.n117 5.56245
R573 w_833_2071.t81 w_833_2071.n116 5.56245
R574 w_833_2071.t81 w_833_2071.n115 5.56245
R575 w_833_2071.t81 w_833_2071.n114 5.56245
R576 w_833_2071.t81 w_833_2071.n113 5.56245
R577 w_833_2071.t81 w_833_2071.n112 5.56245
R578 w_833_2071.t81 w_833_2071.n111 5.56245
R579 w_833_2071.t81 w_833_2071.n122 5.56245
R580 w_833_2071.t81 w_833_2071.n123 5.56245
R581 w_833_2071.t81 w_833_2071.n174 5.56245
R582 w_833_2071.n143 w_833_2071.t102 5.56245
R583 w_833_2071.n196 w_833_2071.n108 4.72356
R584 w_833_2071.n293 w_833_2071.n53 4.25726
R585 w_833_2071.n267 w_833_2071.t0 3.76226
R586 w_833_2071.t0 w_833_2071.n44 3.76226
R587 w_833_2071.t17 w_833_2071.n32 3.76226
R588 w_833_2071.n206 w_833_2071.n56 3.30365
R589 w_833_2071.n208 w_833_2071.n56 3.30365
R590 w_833_2071.n210 w_833_2071.n56 3.30365
R591 w_833_2071.n203 w_833_2071.n56 3.30365
R592 w_833_2071.n201 w_833_2071.n56 3.30365
R593 w_833_2071.n197 w_833_2071.n56 3.30365
R594 w_833_2071.n223 w_833_2071.n54 3.30365
R595 w_833_2071.n225 w_833_2071.n54 3.30365
R596 w_833_2071.n227 w_833_2071.n54 3.30365
R597 w_833_2071.n220 w_833_2071.n54 3.30365
R598 w_833_2071.n218 w_833_2071.n54 3.30365
R599 w_833_2071.n214 w_833_2071.n54 3.30365
R600 w_833_2071.n240 w_833_2071.n57 3.30365
R601 w_833_2071.n242 w_833_2071.n57 3.30365
R602 w_833_2071.n244 w_833_2071.n57 3.30365
R603 w_833_2071.n237 w_833_2071.n57 3.30365
R604 w_833_2071.n235 w_833_2071.n57 3.30365
R605 w_833_2071.n231 w_833_2071.n57 3.30365
R606 w_833_2071.n327 w_833_2071.n20 3.30365
R607 w_833_2071.n327 w_833_2071.n37 3.30365
R608 w_833_2071.n327 w_833_2071.n14 3.30365
R609 w_833_2071.n328 w_833_2071.n327 3.30365
R610 w_833_2071.n327 w_833_2071.n0 3.30365
R611 w_833_2071.n327 w_833_2071.n52 3.30365
R612 w_833_2071.n199 w_833_2071.n56 2.71714
R613 w_833_2071.n216 w_833_2071.n54 2.71714
R614 w_833_2071.n233 w_833_2071.n57 2.71714
R615 w_833_2071.n327 w_833_2071.n5 2.71714
R616 w_833_2071.n204 w_833_2071.n56 2.71618
R617 w_833_2071.n221 w_833_2071.n54 2.71618
R618 w_833_2071.n238 w_833_2071.n57 2.71618
R619 w_833_2071.n327 w_833_2071.n29 2.71618
R620 w_833_2071.n176 w_833_2071.n108 2.10491
R621 w_833_2071.n140 w_833_2071.n108 2.10491
R622 w_833_2071.n264 w_833_2071.n74 1.14089
R623 w_833_2071.n296 w_833_2071.n294 1.13323
R624 w_833_2071.n294 w_833_2071.n252 1.05833
R625 w_833_2071.n264 w_833_2071.n252 1.04625
R626 w_833_2071.n251 w_833_2071.n249 0.80919
R627 w_833_2071.n174 w_833_2071.n173 0.80612
R628 w_833_2071.n144 w_833_2071.n143 0.805774
R629 w_833_2071.n230 w_833_2071.n213 0.794017
R630 w_833_2071.n249 w_833_2071.n247 0.789466
R631 w_833_2071.n247 w_833_2071.n230 0.789466
R632 w_833_2071.n324 w_833_2071.n323 0.722964
R633 w_833_2071.n295 w_833_2071.n66 0.693971
R634 w_833_2071.n213 w_833_2071.n196 0.693879
R635 w_833_2071.n107 w_833_2071.n106 0.6055
R636 w_833_2071.n169 w_833_2071.n168 0.6055
R637 w_833_2071.n177 w_833_2071.n174 0.596545
R638 w_833_2071.n143 w_833_2071.n142 0.569391
R639 w_833_2071.n321 w_833_2071.n101 0.562058
R640 w_833_2071.n75 w_833_2071.n73 0.562058
R641 w_833_2071.n185 w_833_2071.n114 0.562058
R642 w_833_2071.n187 w_833_2071.n113 0.562058
R643 w_833_2071.n189 w_833_2071.n112 0.562058
R644 w_833_2071.n191 w_833_2071.n111 0.562058
R645 w_833_2071.n181 w_833_2071.n122 0.562058
R646 w_833_2071.n179 w_833_2071.n123 0.562058
R647 w_833_2071.n79 w_833_2071.n78 0.561712
R648 w_833_2071.n81 w_833_2071.n80 0.561712
R649 w_833_2071.n83 w_833_2071.n82 0.561712
R650 w_833_2071.n85 w_833_2071.n84 0.561712
R651 w_833_2071.n87 w_833_2071.n86 0.561712
R652 w_833_2071.n89 w_833_2071.n88 0.561712
R653 w_833_2071.n91 w_833_2071.n90 0.561712
R654 w_833_2071.n96 w_833_2071.n95 0.561712
R655 w_833_2071.n98 w_833_2071.n97 0.561712
R656 w_833_2071.n100 w_833_2071.n99 0.561712
R657 w_833_2071.n77 w_833_2071.n76 0.561712
R658 w_833_2071.n137 w_833_2071.n121 0.561712
R659 w_833_2071.n135 w_833_2071.n120 0.561712
R660 w_833_2071.n133 w_833_2071.n119 0.561712
R661 w_833_2071.n131 w_833_2071.n118 0.561712
R662 w_833_2071.n129 w_833_2071.n117 0.561712
R663 w_833_2071.n127 w_833_2071.n116 0.561712
R664 w_833_2071.n125 w_833_2071.n115 0.561712
R665 w_833_2071.n323 w_833_2071.n74 0.50362
R666 w_833_2071.n298 w_833_2071.n79 0.50362
R667 w_833_2071.n300 w_833_2071.n81 0.50362
R668 w_833_2071.n302 w_833_2071.n83 0.50362
R669 w_833_2071.n304 w_833_2071.n85 0.50362
R670 w_833_2071.n306 w_833_2071.n87 0.50362
R671 w_833_2071.n308 w_833_2071.n89 0.50362
R672 w_833_2071.n310 w_833_2071.n91 0.50362
R673 w_833_2071.n314 w_833_2071.n96 0.50362
R674 w_833_2071.n316 w_833_2071.n98 0.50362
R675 w_833_2071.n318 w_833_2071.n100 0.50362
R676 w_833_2071.n105 w_833_2071.n77 0.50362
R677 w_833_2071.n296 w_833_2071.n295 0.50362
R678 w_833_2071.n145 w_833_2071.n121 0.50362
R679 w_833_2071.n147 w_833_2071.n120 0.50362
R680 w_833_2071.n149 w_833_2071.n119 0.50362
R681 w_833_2071.n151 w_833_2071.n118 0.50362
R682 w_833_2071.n153 w_833_2071.n117 0.50362
R683 w_833_2071.n155 w_833_2071.n116 0.50362
R684 w_833_2071.n157 w_833_2071.n115 0.50362
R685 w_833_2071.n321 w_833_2071.n320 0.503274
R686 w_833_2071.n103 w_833_2071.n75 0.503274
R687 w_833_2071.n161 w_833_2071.n114 0.503274
R688 w_833_2071.n163 w_833_2071.n113 0.503274
R689 w_833_2071.n165 w_833_2071.n112 0.503274
R690 w_833_2071.n167 w_833_2071.n111 0.503274
R691 w_833_2071.n170 w_833_2071.n122 0.503274
R692 w_833_2071.n172 w_833_2071.n123 0.503274
R693 w_833_2071.n293 w_833_2071.n264 0.499574
R694 w_833_2071.n294 w_833_2071.n293 0.498883
R695 w_833_2071.n246 w_833_2071.n245 0.37848
R696 w_833_2071.n229 w_833_2071.n228 0.37848
R697 w_833_2071.n212 w_833_2071.n211 0.37848
R698 w_833_2071.n248 w_833_2071.n1 0.37848
R699 w_833_2071.n240 w_833_2071.n239 0.365272
R700 w_833_2071.n223 w_833_2071.n222 0.365272
R701 w_833_2071.n206 w_833_2071.n205 0.365272
R702 w_833_2071.n28 w_833_2071.n20 0.365272
R703 w_833_2071.n235 w_833_2071.n234 0.364033
R704 w_833_2071.n218 w_833_2071.n217 0.364033
R705 w_833_2071.n201 w_833_2071.n200 0.364033
R706 w_833_2071.n4 w_833_2071.n0 0.364033
R707 w_833_2071.n232 w_833_2071.n231 0.357939
R708 w_833_2071.n215 w_833_2071.n214 0.357939
R709 w_833_2071.n198 w_833_2071.n197 0.357939
R710 w_833_2071.n52 w_833_2071.n51 0.357939
R711 w_833_2071.n159 w_833_2071.n109 0.354712
R712 w_833_2071.n242 w_833_2071.n241 0.343272
R713 w_833_2071.n225 w_833_2071.n224 0.343272
R714 w_833_2071.n208 w_833_2071.n207 0.343272
R715 w_833_2071.n37 w_833_2071.n35 0.343272
R716 w_833_2071.n237 w_833_2071.n236 0.342033
R717 w_833_2071.n220 w_833_2071.n219 0.342033
R718 w_833_2071.n203 w_833_2071.n202 0.342033
R719 w_833_2071.n329 w_833_2071.n328 0.342033
R720 w_833_2071.n312 w_833_2071.n92 0.340978
R721 w_833_2071.n244 w_833_2071.n243 0.321272
R722 w_833_2071.n227 w_833_2071.n226 0.321272
R723 w_833_2071.n210 w_833_2071.n209 0.321272
R724 w_833_2071.n36 w_833_2071.n14 0.321272
R725 w_833_2071.n233 w_833_2071.n232 0.320626
R726 w_833_2071.n216 w_833_2071.n215 0.320626
R727 w_833_2071.n199 w_833_2071.n198 0.320626
R728 w_833_2071.n51 w_833_2071.n5 0.320626
R729 w_833_2071.n245 w_833_2071.n244 0.320033
R730 w_833_2071.n228 w_833_2071.n227 0.320033
R731 w_833_2071.n211 w_833_2071.n210 0.320033
R732 w_833_2071.n14 w_833_2071.n1 0.320033
R733 w_833_2071.n239 w_833_2071.n238 0.319212
R734 w_833_2071.n222 w_833_2071.n221 0.319212
R735 w_833_2071.n205 w_833_2071.n204 0.319212
R736 w_833_2071.n29 w_833_2071.n28 0.319212
R737 w_833_2071.n234 w_833_2071.n233 0.315027
R738 w_833_2071.n217 w_833_2071.n216 0.315027
R739 w_833_2071.n200 w_833_2071.n199 0.315027
R740 w_833_2071.n5 w_833_2071.n4 0.315027
R741 w_833_2071.n94 w_833_2071.n93 0.305134
R742 w_833_2071.n102 w_833_2071.n74 0.303
R743 w_833_2071.n103 w_833_2071.n102 0.303
R744 w_833_2071.n104 w_833_2071.n103 0.303
R745 w_833_2071.n105 w_833_2071.n104 0.303
R746 w_833_2071.n106 w_833_2071.n105 0.303
R747 w_833_2071.n320 w_833_2071.n107 0.303
R748 w_833_2071.n320 w_833_2071.n319 0.303
R749 w_833_2071.n319 w_833_2071.n318 0.303
R750 w_833_2071.n318 w_833_2071.n317 0.303
R751 w_833_2071.n317 w_833_2071.n316 0.303
R752 w_833_2071.n316 w_833_2071.n315 0.303
R753 w_833_2071.n315 w_833_2071.n314 0.303
R754 w_833_2071.n314 w_833_2071.n313 0.303
R755 w_833_2071.n313 w_833_2071.n312 0.303
R756 w_833_2071.n312 w_833_2071.n311 0.303
R757 w_833_2071.n311 w_833_2071.n310 0.303
R758 w_833_2071.n310 w_833_2071.n309 0.303
R759 w_833_2071.n309 w_833_2071.n308 0.303
R760 w_833_2071.n308 w_833_2071.n307 0.303
R761 w_833_2071.n307 w_833_2071.n306 0.303
R762 w_833_2071.n306 w_833_2071.n305 0.303
R763 w_833_2071.n305 w_833_2071.n304 0.303
R764 w_833_2071.n304 w_833_2071.n303 0.303
R765 w_833_2071.n303 w_833_2071.n302 0.303
R766 w_833_2071.n302 w_833_2071.n301 0.303
R767 w_833_2071.n301 w_833_2071.n300 0.303
R768 w_833_2071.n300 w_833_2071.n299 0.303
R769 w_833_2071.n299 w_833_2071.n298 0.303
R770 w_833_2071.n298 w_833_2071.n297 0.303
R771 w_833_2071.n297 w_833_2071.n296 0.303
R772 w_833_2071.n173 w_833_2071.n172 0.303
R773 w_833_2071.n172 w_833_2071.n171 0.303
R774 w_833_2071.n171 w_833_2071.n170 0.303
R775 w_833_2071.n170 w_833_2071.n169 0.303
R776 w_833_2071.n168 w_833_2071.n167 0.303
R777 w_833_2071.n167 w_833_2071.n166 0.303
R778 w_833_2071.n166 w_833_2071.n165 0.303
R779 w_833_2071.n165 w_833_2071.n164 0.303
R780 w_833_2071.n164 w_833_2071.n163 0.303
R781 w_833_2071.n163 w_833_2071.n162 0.303
R782 w_833_2071.n162 w_833_2071.n161 0.303
R783 w_833_2071.n161 w_833_2071.n160 0.303
R784 w_833_2071.n160 w_833_2071.n159 0.303
R785 w_833_2071.n159 w_833_2071.n158 0.303
R786 w_833_2071.n158 w_833_2071.n157 0.303
R787 w_833_2071.n157 w_833_2071.n156 0.303
R788 w_833_2071.n156 w_833_2071.n155 0.303
R789 w_833_2071.n155 w_833_2071.n154 0.303
R790 w_833_2071.n154 w_833_2071.n153 0.303
R791 w_833_2071.n153 w_833_2071.n152 0.303
R792 w_833_2071.n152 w_833_2071.n151 0.303
R793 w_833_2071.n151 w_833_2071.n150 0.303
R794 w_833_2071.n150 w_833_2071.n149 0.303
R795 w_833_2071.n149 w_833_2071.n148 0.303
R796 w_833_2071.n148 w_833_2071.n147 0.303
R797 w_833_2071.n147 w_833_2071.n146 0.303
R798 w_833_2071.n146 w_833_2071.n145 0.303
R799 w_833_2071.n145 w_833_2071.n144 0.303
R800 w_833_2071.n245 w_833_2071.n237 0.299272
R801 w_833_2071.n228 w_833_2071.n220 0.299272
R802 w_833_2071.n211 w_833_2071.n203 0.299272
R803 w_833_2071.n328 w_833_2071.n1 0.299272
R804 w_833_2071.n243 w_833_2071.n242 0.298033
R805 w_833_2071.n226 w_833_2071.n225 0.298033
R806 w_833_2071.n209 w_833_2071.n208 0.298033
R807 w_833_2071.n37 w_833_2071.n36 0.298033
R808 w_833_2071.n194 w_833_2071.n110 0.277397
R809 w_833_2071.n236 w_833_2071.n235 0.277272
R810 w_833_2071.n219 w_833_2071.n218 0.277272
R811 w_833_2071.n202 w_833_2071.n201 0.277272
R812 w_833_2071.n329 w_833_2071.n0 0.277272
R813 w_833_2071.n241 w_833_2071.n240 0.276033
R814 w_833_2071.n224 w_833_2071.n223 0.276033
R815 w_833_2071.n207 w_833_2071.n206 0.276033
R816 w_833_2071.n35 w_833_2071.n20 0.276033
R817 w_833_2071.n88 w_833_2071.n63 0.198759
R818 w_833_2071.n127 w_833_2071.n126 0.198419
R819 w_833_2071.n193 w_833_2071.n192 0.191425
R820 w_833_2071.n322 w_833_2071.n72 0.191086
R821 w_833_2071.n78 w_833_2071.n66 0.191086
R822 w_833_2071.n90 w_833_2071.n62 0.187772
R823 w_833_2071.n125 w_833_2071.n124 0.187772
R824 w_833_2071.n78 w_833_2071.n67 0.186494
R825 w_833_2071.n137 w_833_2071.n136 0.186494
R826 w_833_2071.n322 w_833_2071.n59 0.184092
R827 w_833_2071.n193 w_833_2071.n182 0.183752
R828 w_833_2071.n101 w_833_2071.n60 0.180439
R829 w_833_2071.n80 w_833_2071.n68 0.180439
R830 w_833_2071.n191 w_833_2071.n190 0.180439
R831 w_833_2071.n135 w_833_2071.n134 0.180439
R832 w_833_2071.n93 w_833_2071.n70 0.176759
R833 w_833_2071.n88 w_833_2071.n69 0.176419
R834 w_833_2071.n128 w_833_2071.n127 0.176419
R835 w_833_2071.n76 w_833_2071.n58 0.173106
R836 w_833_2071.n181 w_833_2071.n180 0.173106
R837 w_833_2071.n184 w_833_2071.n183 0.172752
R838 w_833_2071.n82 w_833_2071.n65 0.169425
R839 w_833_2071.n189 w_833_2071.n188 0.169425
R840 w_833_2071.n99 w_833_2071.n61 0.169086
R841 w_833_2071.n133 w_833_2071.n132 0.169086
R842 w_833_2071.n95 w_833_2071.n71 0.165772
R843 w_833_2071.n86 w_833_2071.n64 0.165772
R844 w_833_2071.n186 w_833_2071.n185 0.165772
R845 w_833_2071.n130 w_833_2071.n129 0.165772
R846 w_833_2071.n324 w_833_2071.n73 0.162092
R847 w_833_2071.n179 w_833_2071.n178 0.161752
R848 w_833_2071.n97 w_833_2071.n71 0.158439
R849 w_833_2071.n84 w_833_2071.n64 0.158439
R850 w_833_2071.n187 w_833_2071.n186 0.158439
R851 w_833_2071.n131 w_833_2071.n130 0.158439
R852 w_833_2071.n97 w_833_2071.n61 0.154759
R853 w_833_2071.n132 w_833_2071.n131 0.154759
R854 w_833_2071.n84 w_833_2071.n65 0.154419
R855 w_833_2071.n188 w_833_2071.n187 0.154419
R856 w_833_2071.n141 w_833_2071.n138 0.152939
R857 w_833_2071.n73 w_833_2071.n58 0.151106
R858 w_833_2071.n180 w_833_2071.n179 0.151106
R859 w_833_2071.n86 w_833_2071.n69 0.147425
R860 w_833_2071.n185 w_833_2071.n184 0.147425
R861 w_833_2071.n129 w_833_2071.n128 0.147425
R862 w_833_2071.n95 w_833_2071.n70 0.147086
R863 w_833_2071.n195 w_833_2071.n109 0.146921
R864 w_833_2071.n99 w_833_2071.n60 0.143772
R865 w_833_2071.n82 w_833_2071.n68 0.143772
R866 w_833_2071.n190 w_833_2071.n189 0.143772
R867 w_833_2071.n134 w_833_2071.n133 0.143772
R868 w_833_2071.n182 w_833_2071.n181 0.140092
R869 w_833_2071.n76 w_833_2071.n59 0.139752
R870 w_833_2071.n80 w_833_2071.n67 0.137241
R871 w_833_2071.n136 w_833_2071.n135 0.137241
R872 w_833_2071.n93 w_833_2071.n62 0.136439
R873 w_833_2071.n124 w_833_2071.n110 0.136439
R874 w_833_2071.n101 w_833_2071.n72 0.132759
R875 w_833_2071.n192 w_833_2071.n191 0.132419
R876 w_833_2071.n138 w_833_2071.n137 0.129106
R877 w_833_2071.n178 w_833_2071.n177 0.127259
R878 w_833_2071.n126 w_833_2071.n125 0.125425
R879 w_833_2071.n90 w_833_2071.n63 0.125086
R880 w_833_2071.n250 w_833_2071.n94 0.1105
R881 w_833_2071.n250 w_833_2071.n92 0.0990487
R882 w_833_2071.n195 w_833_2071.n194 0.0763621
R883 w_833_2071.n142 w_833_2071.n141 0.0353333
R884 w_833_2071.n183 w_833_2071.n110 0.00416667
R885 vinp.n0 vinp.t16 15.8289
R886 vinp.n22 vinp.t27 15.8289
R887 vinp.n15 vinp.t21 15.6055
R888 vinp.n7 vinp.t12 15.6055
R889 vinp.n6 vinp.t13 15.2239
R890 vinp.n5 vinp.t18 15.2239
R891 vinp.n4 vinp.t24 15.2239
R892 vinp.n3 vinp.t7 15.2239
R893 vinp.n2 vinp.t5 15.2239
R894 vinp.n1 vinp.t14 15.2239
R895 vinp.n0 vinp.t9 15.2239
R896 vinp.n28 vinp.t26 15.2239
R897 vinp.n27 vinp.t31 15.2239
R898 vinp.n26 vinp.t2 15.2239
R899 vinp.n25 vinp.t15 15.2239
R900 vinp.n24 vinp.t10 15.2239
R901 vinp.n23 vinp.t25 15.2239
R902 vinp.n22 vinp.t19 15.2239
R903 vinp.n15 vinp.t28 15.0005
R904 vinp.n16 vinp.t8 15.0005
R905 vinp.n17 vinp.t1 15.0005
R906 vinp.n18 vinp.t4 15.0005
R907 vinp.n19 vinp.t0 15.0005
R908 vinp.n20 vinp.t3 15.0005
R909 vinp.n21 vinp.t20 15.0005
R910 vinp.n7 vinp.t17 15.0005
R911 vinp.n8 vinp.t6 15.0005
R912 vinp.n9 vinp.t23 15.0005
R913 vinp.n10 vinp.t30 15.0005
R914 vinp.n11 vinp.t22 15.0005
R915 vinp.n12 vinp.t29 15.0005
R916 vinp.n13 vinp.t11 15.0005
R917 vinp vinp.n30 12.0616
R918 vinp.n14 vinp 10.4452
R919 vinp.n29 vinp 10.1782
R920 vinp.n29 vinp 9.53331
R921 vinp.n14 vinp 9.26175
R922 vinp vinp.n6 4.90238
R923 vinp vinp.n28 4.90238
R924 vinp.n1 vinp.n0 0.6055
R925 vinp.n2 vinp.n1 0.6055
R926 vinp.n3 vinp.n2 0.6055
R927 vinp.n4 vinp.n3 0.6055
R928 vinp.n5 vinp.n4 0.6055
R929 vinp.n6 vinp.n5 0.6055
R930 vinp.n23 vinp.n22 0.6055
R931 vinp.n24 vinp.n23 0.6055
R932 vinp.n25 vinp.n24 0.6055
R933 vinp.n26 vinp.n25 0.6055
R934 vinp.n27 vinp.n26 0.6055
R935 vinp.n28 vinp.n27 0.6055
R936 vinp.n16 vinp.n15 0.6055
R937 vinp.n17 vinp.n16 0.6055
R938 vinp.n18 vinp.n17 0.6055
R939 vinp.n19 vinp.n18 0.6055
R940 vinp.n20 vinp.n19 0.6055
R941 vinp.n21 vinp.n20 0.6055
R942 vinp.n8 vinp.n7 0.6055
R943 vinp.n9 vinp.n8 0.6055
R944 vinp.n10 vinp.n9 0.6055
R945 vinp.n11 vinp.n10 0.6055
R946 vinp.n12 vinp.n11 0.6055
R947 vinp.n13 vinp.n12 0.6055
R948 vinp.n30 vinp.n29 0.425328
R949 vinp vinp.n21 0.333938
R950 vinp vinp.n13 0.333938
R951 vinp.n30 vinp.n14 0.241741
R952 a_610_6649.n28 a_610_6649.t10 18.8663
R953 a_610_6649.n0 a_610_6649.t3 18.8633
R954 a_610_6649.n32 a_610_6649.t4 18.619
R955 a_610_6649.n24 a_610_6649.t11 18.619
R956 a_610_6649.n30 a_610_6649.t2 18.1315
R957 a_610_6649.n29 a_610_6649.t1 18.1315
R958 a_610_6649.n28 a_610_6649.t7 18.1315
R959 a_610_6649.n36 a_610_6649.t8 18.1285
R960 a_610_6649.n0 a_610_6649.t14 18.1285
R961 a_610_6649.t15 a_610_6649.n37 18.1285
R962 a_610_6649.n34 a_610_6649.t0 17.8842
R963 a_610_6649.n33 a_610_6649.t12 17.8842
R964 a_610_6649.n32 a_610_6649.t5 17.8842
R965 a_610_6649.n26 a_610_6649.t9 17.8842
R966 a_610_6649.n25 a_610_6649.t6 17.8842
R967 a_610_6649.n24 a_610_6649.t13 17.8842
R968 a_610_6649.n27 a_610_6649.n23 15.7467
R969 a_610_6649.n35 a_610_6649.n34 13.4687
R970 a_610_6649.n27 a_610_6649.n26 13.4687
R971 a_610_6649.n36 a_610_6649.n35 11.1279
R972 a_610_6649.n23 a_610_6649.n1 10.8121
R973 a_610_6649.n31 a_610_6649.n30 10.3711
R974 a_610_6649.n23 a_610_6649.n22 9.36767
R975 a_610_6649.n2 a_610_6649.t23 5.63764
R976 a_610_6649.n11 a_610_6649.t21 5.63764
R977 a_610_6649.n21 a_610_6649.t17 5.63764
R978 a_610_6649.n14 a_610_6649.t19 5.63764
R979 a_610_6649.n2 a_610_6649.n1 5.47498
R980 a_610_6649.n22 a_610_6649.n11 5.47498
R981 a_610_6649.n22 a_610_6649.n21 4.57374
R982 a_610_6649.n14 a_610_6649.n1 4.57374
R983 a_610_6649.n8 a_610_6649.t34 4.42794
R984 a_610_6649.n3 a_610_6649.t28 4.42666
R985 a_610_6649.n12 a_610_6649.t29 4.42666
R986 a_610_6649.n18 a_610_6649.t35 4.42557
R987 a_610_6649.n3 a_610_6649.t32 2.82253
R988 a_610_6649.n4 a_610_6649.t26 2.82253
R989 a_610_6649.n6 a_610_6649.t22 2.82253
R990 a_610_6649.n7 a_610_6649.t27 2.82253
R991 a_610_6649.n9 a_610_6649.t20 2.82253
R992 a_610_6649.n8 a_610_6649.t30 2.82253
R993 a_610_6649.n12 a_610_6649.t33 2.82253
R994 a_610_6649.n13 a_610_6649.t24 2.82253
R995 a_610_6649.n16 a_610_6649.t18 2.82253
R996 a_610_6649.n17 a_610_6649.t25 2.82253
R997 a_610_6649.n19 a_610_6649.t16 2.82253
R998 a_610_6649.n18 a_610_6649.t31 2.82253
R999 a_610_6649.n4 a_610_6649.n3 1.60563
R1000 a_610_6649.n7 a_610_6649.n6 1.60563
R1001 a_610_6649.n9 a_610_6649.n8 1.60563
R1002 a_610_6649.n13 a_610_6649.n12 1.60563
R1003 a_610_6649.n17 a_610_6649.n16 1.60563
R1004 a_610_6649.n19 a_610_6649.n18 1.60563
R1005 a_610_6649.n35 a_610_6649.n31 1.4635
R1006 a_610_6649.n5 a_610_6649.n4 0.803704
R1007 a_610_6649.n10 a_610_6649.n7 0.803704
R1008 a_610_6649.n15 a_610_6649.n13 0.803704
R1009 a_610_6649.n20 a_610_6649.n17 0.803704
R1010 a_610_6649.n6 a_610_6649.n5 0.802423
R1011 a_610_6649.n10 a_610_6649.n9 0.802423
R1012 a_610_6649.n16 a_610_6649.n15 0.802423
R1013 a_610_6649.n20 a_610_6649.n19 0.802423
R1014 a_610_6649.n31 a_610_6649.n27 0.7463
R1015 a_610_6649.n33 a_610_6649.n32 0.7353
R1016 a_610_6649.n34 a_610_6649.n33 0.7353
R1017 a_610_6649.n29 a_610_6649.n28 0.7353
R1018 a_610_6649.n30 a_610_6649.n29 0.7353
R1019 a_610_6649.n25 a_610_6649.n24 0.7353
R1020 a_610_6649.n26 a_610_6649.n25 0.7353
R1021 a_610_6649.n37 a_610_6649.n36 0.7353
R1022 a_610_6649.n37 a_610_6649.n0 0.7353
R1023 a_610_6649.n5 a_610_6649.n2 0.390831
R1024 a_610_6649.n11 a_610_6649.n10 0.390831
R1025 a_610_6649.n21 a_610_6649.n20 0.390831
R1026 a_610_6649.n15 a_610_6649.n14 0.390831
R1027 vinn.n15 vinn.t28 15.8289
R1028 vinn.n7 vinn.t18 15.8289
R1029 vinn.n0 vinn.t9 15.6055
R1030 vinn.n22 vinn.t20 15.6055
R1031 vinn.n21 vinn.t26 15.2239
R1032 vinn.n20 vinn.t0 15.2239
R1033 vinn.n19 vinn.t4 15.2239
R1034 vinn.n18 vinn.t13 15.2239
R1035 vinn.n17 vinn.t10 15.2239
R1036 vinn.n16 vinn.t27 15.2239
R1037 vinn.n15 vinn.t21 15.2239
R1038 vinn.n13 vinn.t15 15.2239
R1039 vinn.n12 vinn.t22 15.2239
R1040 vinn.n11 vinn.t29 15.2239
R1041 vinn.n10 vinn.t8 15.2239
R1042 vinn.n9 vinn.t5 15.2239
R1043 vinn.n8 vinn.t14 15.2239
R1044 vinn.n7 vinn.t12 15.2239
R1045 vinn.n0 vinn.t11 15.0005
R1046 vinn.n1 vinn.t2 15.0005
R1047 vinn.n2 vinn.t19 15.0005
R1048 vinn.n3 vinn.t24 15.0005
R1049 vinn.n4 vinn.t16 15.0005
R1050 vinn.n5 vinn.t23 15.0005
R1051 vinn.n6 vinn.t7 15.0005
R1052 vinn.n22 vinn.t25 15.0005
R1053 vinn.n23 vinn.t6 15.0005
R1054 vinn.n24 vinn.t31 15.0005
R1055 vinn.n25 vinn.t3 15.0005
R1056 vinn.n26 vinn.t30 15.0005
R1057 vinn.n27 vinn.t1 15.0005
R1058 vinn.n28 vinn.t17 15.0005
R1059 vinn vinn.n30 11.8039
R1060 vinn.n29 vinn 10.6252
R1061 vinn.n14 vinn 10.3506
R1062 vinn.n14 vinn 9.95612
R1063 vinn.n29 vinn 9.68456
R1064 vinn vinn.n21 4.90238
R1065 vinn vinn.n13 4.90238
R1066 vinn.n1 vinn.n0 0.6055
R1067 vinn.n2 vinn.n1 0.6055
R1068 vinn.n3 vinn.n2 0.6055
R1069 vinn.n4 vinn.n3 0.6055
R1070 vinn.n5 vinn.n4 0.6055
R1071 vinn.n6 vinn.n5 0.6055
R1072 vinn.n23 vinn.n22 0.6055
R1073 vinn.n24 vinn.n23 0.6055
R1074 vinn.n25 vinn.n24 0.6055
R1075 vinn.n26 vinn.n25 0.6055
R1076 vinn.n27 vinn.n26 0.6055
R1077 vinn.n28 vinn.n27 0.6055
R1078 vinn.n16 vinn.n15 0.6055
R1079 vinn.n17 vinn.n16 0.6055
R1080 vinn.n18 vinn.n17 0.6055
R1081 vinn.n19 vinn.n18 0.6055
R1082 vinn.n20 vinn.n19 0.6055
R1083 vinn.n21 vinn.n20 0.6055
R1084 vinn.n8 vinn.n7 0.6055
R1085 vinn.n9 vinn.n8 0.6055
R1086 vinn.n10 vinn.n9 0.6055
R1087 vinn.n11 vinn.n10 0.6055
R1088 vinn.n12 vinn.n11 0.6055
R1089 vinn.n13 vinn.n12 0.6055
R1090 vinn.n30 vinn.n14 0.548224
R1091 vinn.n30 vinn.n29 0.364638
R1092 vinn vinn.n6 0.333938
R1093 vinn vinn.n28 0.333938
R1094 vout.n15 vout.t12 18.8648
R1095 vout.n7 vout.t16 18.8648
R1096 vout.n11 vout.t13 18.6205
R1097 vout.n4 vout.t9 18.6175
R1098 vout.n17 vout.t19 18.13
R1099 vout.n16 vout.t14 18.13
R1100 vout.n15 vout.t11 18.13
R1101 vout.n9 vout.t10 18.13
R1102 vout.n8 vout.t4 18.13
R1103 vout.n7 vout.t5 18.13
R1104 vout.n13 vout.t15 17.8857
R1105 vout.n12 vout.t17 17.8857
R1106 vout.n11 vout.t6 17.8857
R1107 vout.n6 vout.t7 17.8827
R1108 vout.n5 vout.t8 17.8827
R1109 vout.n4 vout.t18 17.8827
R1110 vout.n3 vout.n2 15.106
R1111 vout.n2 vout.n0 13.7009
R1112 vout.n18 vout.n17 13.4665
R1113 vout.n10 vout.n9 13.4665
R1114 vout.n10 vout.n6 11.8385
R1115 vout.n0 vout.t0 11.1117
R1116 vout.n1 vout.t2 11.1117
R1117 vout.n3 vout 10.8815
R1118 vout.n14 vout.n13 10.3689
R1119 vout.n0 vout.t1 10.2104
R1120 vout.n1 vout.t3 10.2104
R1121 vout.n2 vout.n1 9.36767
R1122 vout.n18 vout.n14 1.4591
R1123 vout vout.n3 0.8673
R1124 vout.n14 vout.n10 0.7507
R1125 vout.n16 vout.n15 0.7353
R1126 vout.n17 vout.n16 0.7353
R1127 vout.n12 vout.n11 0.7353
R1128 vout.n13 vout.n12 0.7353
R1129 vout.n8 vout.n7 0.7353
R1130 vout.n9 vout.n8 0.7353
R1131 vout.n5 vout.n4 0.7353
R1132 vout.n6 vout.n5 0.7353
R1133 vout vout.n18 0.3041
C0 vinp vout 0.91461f
C1 vinn vout 2.65413f
C2 vinp vdda 0.13084f
C3 vinn vdda 0.43281f
C4 vinn vinp 6.92099f
C5 vdda vout 1.75926f
C6 w_609_1847# vdda 0.26354f
C7 ibias vssa 20.1072f
C8 vinp vssa 5.42415f
C9 vinn vssa 5.82446f
C10 vout vssa 2.67846f
C11 vdda vssa 5.61529f
C12 w_609_1847# vssa 0.11231f $ **FLOATING
C13 vout.t0 vssa 0.19789f
C14 vout.t1 vssa 0.1781f
C15 vout.n0 vssa 0.82078f
C16 vout.t2 vssa 0.19789f
C17 vout.t3 vssa 0.17811f
C18 vout.n1 vssa 0.57261f
C19 vout.n2 vssa 1.72598f
C20 vout.n3 vssa 0.89068f
C21 vout.t9 vssa 0.30436f
C22 vout.t18 vssa 0.32571f
C23 vout.n4 vssa -0.24134f
C24 vout.t8 vssa 0.32571f
C25 vout.n5 vssa 0.27814f
C26 vout.t7 vssa 0.32571f
C27 vout.n6 vssa 0.46652f
C28 vout.t16 vssa 0.33846f
C29 vout.t5 vssa 0.33883f
C30 vout.n7 vssa 0.27948f
C31 vout.t4 vssa 0.33883f
C32 vout.n8 vssa 0.28863f
C33 vout.t10 vssa 0.33883f
C34 vout.n9 vssa 0.86464f
C35 vout.n10 vssa 0.47736f
C36 vout.t13 vssa 0.30438f
C37 vout.t6 vssa 0.32572f
C38 vout.n11 vssa -0.24136f
C39 vout.t17 vssa 0.32572f
C40 vout.n12 vssa 0.27814f
C41 vout.t15 vssa 0.32572f
C42 vout.n13 vssa 0.44606f
C43 vout.n14 vssa 0.21944f
C44 vout.t12 vssa 0.33846f
C45 vout.t11 vssa 0.33883f
C46 vout.n15 vssa 0.27948f
C47 vout.t14 vssa 0.33883f
C48 vout.n16 vssa 0.28863f
C49 vout.t19 vssa 0.33883f
C50 vout.n17 vssa 0.86464f
C51 vout.n18 vssa 0.29405f
C52 vinn.t9 vssa 0.43961f
C53 vinn.t11 vssa 0.43721f
C54 vinn.n0 vssa 0.15546f
C55 vinn.t2 vssa 0.43721f
C56 vinn.t19 vssa 0.43721f
C57 vinn.t24 vssa 0.43721f
C58 vinn.t16 vssa 0.43721f
C59 vinn.t23 vssa 0.43721f
C60 vinn.t7 vssa 0.43721f
C61 vinn.t15 vssa 0.43767f
C62 vinn.t22 vssa 0.43767f
C63 vinn.t29 vssa 0.43767f
C64 vinn.t8 vssa 0.43767f
C65 vinn.t5 vssa 0.43767f
C66 vinn.t14 vssa 0.43767f
C67 vinn.t12 vssa 0.43767f
C68 vinn.t18 vssa 0.44171f
C69 vinn.n7 vssa 0.24653f
C70 vinn.n8 vssa 0.14488f
C71 vinn.n9 vssa 0.14488f
C72 vinn.n10 vssa 0.14488f
C73 vinn.n11 vssa 0.14488f
C74 vinn.n12 vssa 0.14488f
C75 vinn.n13 vssa 0.48512f
C76 vinn.n14 vssa 0.64269f
C77 vinn.t26 vssa 0.43767f
C78 vinn.t0 vssa 0.43767f
C79 vinn.t4 vssa 0.43767f
C80 vinn.t13 vssa 0.43767f
C81 vinn.t10 vssa 0.43767f
C82 vinn.t27 vssa 0.43767f
C83 vinn.t21 vssa 0.43767f
C84 vinn.t28 vssa 0.44171f
C85 vinn.n15 vssa 0.24653f
C86 vinn.n16 vssa 0.14488f
C87 vinn.n17 vssa 0.14488f
C88 vinn.n18 vssa 0.14488f
C89 vinn.n19 vssa 0.14488f
C90 vinn.n20 vssa 0.14488f
C91 vinn.n21 vssa 0.48512f
C92 vinn.t20 vssa 0.43961f
C93 vinn.t25 vssa 0.43721f
C94 vinn.n22 vssa 0.15546f
C95 vinn.t6 vssa 0.43721f
C96 vinn.t31 vssa 0.43721f
C97 vinn.t3 vssa 0.43721f
C98 vinn.t30 vssa 0.43721f
C99 vinn.t1 vssa 0.43721f
C100 vinn.t17 vssa 0.43721f
C101 vinn.n29 vssa 0.58496f
C102 vinn.n30 vssa 0.42003f
C103 a_610_6649.t3 vssa 0.27916f
C104 a_610_6649.t14 vssa 0.2973f
C105 a_610_6649.n0 vssa -0.19426f
C106 a_610_6649.n1 vssa 0.44276f
C107 a_610_6649.t21 vssa 0.12354f
C108 a_610_6649.t27 vssa 0.84459f
C109 a_610_6649.t22 vssa 0.84459f
C110 a_610_6649.t23 vssa 0.12354f
C111 a_610_6649.t26 vssa 0.84459f
C112 a_610_6649.t32 vssa 0.84459f
C113 a_610_6649.t28 vssa 0.88453f
C114 a_610_6649.n3 vssa 0.19391f
C115 a_610_6649.t34 vssa 0.88353f
C116 a_610_6649.t30 vssa 0.84459f
C117 a_610_6649.n8 vssa 0.19212f
C118 a_610_6649.t20 vssa 0.84459f
C119 a_610_6649.t17 vssa 0.12354f
C120 a_610_6649.t25 vssa 0.84459f
C121 a_610_6649.t18 vssa 0.84459f
C122 a_610_6649.t24 vssa 0.84459f
C123 a_610_6649.t33 vssa 0.84459f
C124 a_610_6649.t29 vssa 0.88453f
C125 a_610_6649.n12 vssa 0.19391f
C126 a_610_6649.t19 vssa 0.12354f
C127 a_610_6649.t35 vssa 0.88352f
C128 a_610_6649.t31 vssa 0.84459f
C129 a_610_6649.n18 vssa 0.19213f
C130 a_610_6649.t16 vssa 0.84459f
C131 a_610_6649.n22 vssa 0.41061f
C132 a_610_6649.n23 vssa 1.16749f
C133 a_610_6649.t11 vssa 0.28535f
C134 a_610_6649.t13 vssa 0.28603f
C135 a_610_6649.n24 vssa 0.22769f
C136 a_610_6649.t6 vssa 0.28603f
C137 a_610_6649.n25 vssa 0.24425f
C138 a_610_6649.t9 vssa 0.28603f
C139 a_610_6649.n26 vssa 0.75033f
C140 a_610_6649.n27 vssa 0.82741f
C141 a_610_6649.t10 vssa 0.27967f
C142 a_610_6649.t7 vssa 0.29779f
C143 a_610_6649.n28 vssa -0.19337f
C144 a_610_6649.t1 vssa 0.29779f
C145 a_610_6649.n29 vssa 0.25369f
C146 a_610_6649.t2 vssa 0.29779f
C147 a_610_6649.n30 vssa 0.40144f
C148 a_610_6649.n31 vssa 0.19275f
C149 a_610_6649.t4 vssa 0.28535f
C150 a_610_6649.t5 vssa 0.28603f
C151 a_610_6649.n32 vssa 0.22769f
C152 a_610_6649.t12 vssa 0.28603f
C153 a_610_6649.n33 vssa 0.24425f
C154 a_610_6649.t0 vssa 0.28603f
C155 a_610_6649.n34 vssa 0.75033f
C156 a_610_6649.n35 vssa 0.32936f
C157 a_610_6649.t8 vssa 0.2973f
C158 a_610_6649.n36 vssa 0.40367f
C159 a_610_6649.n37 vssa 0.25324f
C160 a_610_6649.t15 vssa 0.2973f
C161 vinp.t13 vssa 0.42436f
C162 vinp.t18 vssa 0.42436f
C163 vinp.t24 vssa 0.42436f
C164 vinp.t7 vssa 0.42436f
C165 vinp.t5 vssa 0.42436f
C166 vinp.t14 vssa 0.42436f
C167 vinp.t9 vssa 0.42436f
C168 vinp.t16 vssa 0.42827f
C169 vinp.n0 vssa 0.23903f
C170 vinp.n1 vssa 0.14048f
C171 vinp.n2 vssa 0.14048f
C172 vinp.n3 vssa 0.14048f
C173 vinp.n4 vssa 0.14048f
C174 vinp.n5 vssa 0.14048f
C175 vinp.n6 vssa 0.47036f
C176 vinp.t12 vssa 0.42624f
C177 vinp.t17 vssa 0.4239f
C178 vinp.n7 vssa 0.15074f
C179 vinp.t6 vssa 0.4239f
C180 vinp.t23 vssa 0.4239f
C181 vinp.t30 vssa 0.4239f
C182 vinp.t22 vssa 0.4239f
C183 vinp.t29 vssa 0.4239f
C184 vinp.t11 vssa 0.4239f
C185 vinp.n14 vssa 0.65751f
C186 vinp.t21 vssa 0.42624f
C187 vinp.t28 vssa 0.4239f
C188 vinp.n15 vssa 0.15074f
C189 vinp.t8 vssa 0.4239f
C190 vinp.t1 vssa 0.4239f
C191 vinp.t4 vssa 0.4239f
C192 vinp.t0 vssa 0.4239f
C193 vinp.t3 vssa 0.4239f
C194 vinp.t20 vssa 0.4239f
C195 vinp.t26 vssa 0.42436f
C196 vinp.t31 vssa 0.42436f
C197 vinp.t2 vssa 0.42436f
C198 vinp.t15 vssa 0.42436f
C199 vinp.t10 vssa 0.42436f
C200 vinp.t25 vssa 0.42436f
C201 vinp.t19 vssa 0.42436f
C202 vinp.t27 vssa 0.42827f
C203 vinp.n22 vssa 0.23903f
C204 vinp.n23 vssa 0.14048f
C205 vinp.n24 vssa 0.14048f
C206 vinp.n25 vssa 0.14048f
C207 vinp.n26 vssa 0.14048f
C208 vinp.n27 vssa 0.14048f
C209 vinp.n28 vssa 0.47036f
C210 vinp.n29 vssa 0.71753f
C211 vinp.n30 vssa 0.3488f
C212 w_833_2071.t38 vssa 0.38148f
C213 w_833_2071.n2 vssa 0.172f
C214 w_833_2071.n3 vssa 0.24367f
C215 w_833_2071.n6 vssa 0.24367f
C216 w_833_2071.n7 vssa 0.24367f
C217 w_833_2071.n8 vssa 0.11467f
C218 w_833_2071.n9 vssa 0.24367f
C219 w_833_2071.n10 vssa 0.24367f
C220 w_833_2071.n11 vssa 0.24367f
C221 w_833_2071.n13 vssa 0.20067f
C222 w_833_2071.n15 vssa 0.24367f
C223 w_833_2071.n16 vssa 0.24367f
C224 w_833_2071.n17 vssa 0.24367f
C225 w_833_2071.n18 vssa 0.14334f
C226 w_833_2071.n19 vssa 0.24367f
C227 w_833_2071.n21 vssa 0.24367f
C228 w_833_2071.n22 vssa 0.24367f
C229 w_833_2071.n24 vssa 0.215f
C230 w_833_2071.n25 vssa 1.73435f
C231 w_833_2071.n26 vssa 0.24367f
C232 w_833_2071.n27 vssa 0.24367f
C233 w_833_2071.n30 vssa 0.258f
C234 w_833_2071.n31 vssa 0.18634f
C235 w_833_2071.n33 vssa 0.24367f
C236 w_833_2071.n34 vssa 0.24367f
C237 w_833_2071.n38 vssa 0.24367f
C238 w_833_2071.n39 vssa 0.10033f
C239 w_833_2071.n40 vssa 0.24367f
C240 w_833_2071.n41 vssa 0.24367f
C241 w_833_2071.n42 vssa 0.24367f
C242 w_833_2071.n43 vssa 0.15767f
C243 w_833_2071.n44 vssa 0.22934f
C244 w_833_2071.n45 vssa 0.24367f
C245 w_833_2071.n46 vssa 0.24367f
C246 w_833_2071.n47 vssa 0.215f
C247 w_833_2071.n49 vssa 0.24367f
C248 w_833_2071.n50 vssa 0.24367f
C249 w_833_2071.n53 vssa 0.10586f
C250 w_833_2071.n54 vssa 0.38768f
C251 w_833_2071.n55 vssa 0.38768f
C252 w_833_2071.n56 vssa 0.38768f
C253 w_833_2071.n57 vssa 0.38768f
C254 w_833_2071.n108 vssa 0.19108f
C255 w_833_2071.n139 vssa 0.29762f
C256 w_833_2071.n140 vssa 0.13119f
C257 w_833_2071.n175 vssa 0.29736f
C258 w_833_2071.n176 vssa 0.13119f
C259 w_833_2071.t81 vssa 0.54392f
C260 w_833_2071.n251 vssa 0.11784f
C261 w_833_2071.n252 vssa 0.13574f
C262 w_833_2071.t15 vssa 0.215f
C263 w_833_2071.t56 vssa 0.215f
C264 w_833_2071.n254 vssa 0.20067f
C265 w_833_2071.n255 vssa 0.24367f
C266 w_833_2071.n256 vssa 0.24367f
C267 w_833_2071.n257 vssa 0.24367f
C268 w_833_2071.t30 vssa 0.215f
C269 w_833_2071.n258 vssa 0.129f
C270 w_833_2071.n259 vssa 0.24367f
C271 w_833_2071.n260 vssa 0.24367f
C272 w_833_2071.n261 vssa 0.24367f
C273 w_833_2071.t28 vssa 0.215f
C274 w_833_2071.t2 vssa 0.215f
C275 w_833_2071.n263 vssa 0.215f
C276 w_833_2071.n265 vssa 0.24367f
C277 w_833_2071.n266 vssa 0.24367f
C278 w_833_2071.n267 vssa 0.22934f
C279 w_833_2071.t24 vssa 0.215f
C280 w_833_2071.n268 vssa 0.15767f
C281 w_833_2071.n269 vssa 0.24367f
C282 w_833_2071.n270 vssa 0.24367f
C283 w_833_2071.n271 vssa 0.24367f
C284 w_833_2071.t23 vssa 0.215f
C285 w_833_2071.n272 vssa 0.10033f
C286 w_833_2071.n273 vssa 0.24367f
C287 w_833_2071.n274 vssa 0.24367f
C288 w_833_2071.n275 vssa 0.24367f
C289 w_833_2071.t12 vssa 0.215f
C290 w_833_2071.n276 vssa 0.20067f
C291 w_833_2071.t6 vssa 0.215f
C292 w_833_2071.n278 vssa 0.24367f
C293 w_833_2071.n279 vssa 0.24367f
C294 w_833_2071.n280 vssa 0.24367f
C295 w_833_2071.t4 vssa 0.215f
C296 w_833_2071.n281 vssa 0.11467f
C297 w_833_2071.n282 vssa 0.24367f
C298 w_833_2071.n283 vssa 0.24367f
C299 w_833_2071.n284 vssa 0.24367f
C300 w_833_2071.t9 vssa 0.215f
C301 w_833_2071.n285 vssa 0.172f
C302 w_833_2071.t52 vssa 0.24367f
C303 w_833_2071.n286 vssa 0.24367f
C304 w_833_2071.n287 vssa 0.24367f
C305 w_833_2071.t17 vssa 0.215f
C306 w_833_2071.n288 vssa 0.22934f
C307 w_833_2071.t19 vssa 0.215f
C308 w_833_2071.n290 vssa 0.258f
C309 w_833_2071.n291 vssa 0.24367f
C310 w_833_2071.n292 vssa 0.24367f
C311 w_833_2071.n293 vssa 0.93734f
C312 w_833_2071.t75 vssa 0.54392f
C313 w_833_2071.n325 vssa 0.38768f
C314 w_833_2071.n326 vssa 1.48569f
C315 w_833_2071.n327 vssa 0.38768f
.ends

