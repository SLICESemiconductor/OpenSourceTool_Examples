* NGSPICE file created from sg13g2_IOPadIOVss_flat.ext - technology: ihp-sg13g2

.subckt sg13g2_IOPadIOVss_flat iovss vdd vss iovdd
X0 iovss.t4 iovdd.t0 dpantenna l=27.78u w=1.26u
X1 iovss.t5 iovdd.t0 dpantenna l=27.78u w=1.26u
X2 iovss.t3 iovss.t2 dantenna l=27.78u w=1.26u
X3 iovss.t1 iovss.t0 dantenna l=27.78u w=1.26u
R0 iovss.n3104 iovss.n904 21.7649
R1 iovss.n1113 iovss.n1108 9.0005
R2 iovss.n1114 iovss.n1108 9.0005
R3 iovss.n3101 iovss.n1108 9.0005
R4 iovss.n3108 iovss.n3107 9.0005
R5 iovss.n3108 iovss.n1057 9.0005
R6 iovss.n3100 iovss.n1113 9.0005
R7 iovss.n3100 iovss.n1114 9.0005
R8 iovss.n3101 iovss.n3100 9.0005
R9 iovss.n1057 iovss.n965 9.0005
R10 iovss.n3107 iovss.n965 9.0005
R11 iovss.n3077 iovss.n3076 9.0005
R12 iovss.n3076 iovss.n2930 9.0005
R13 iovss.n3078 iovss.n3077 9.0005
R14 iovss.n3078 iovss.n2930 9.0005
R15 iovss.n2093 iovss.n2092 9.0005
R16 iovss.n2089 iovss.n2015 9.0005
R17 iovss.n2089 iovss.n2017 9.0005
R18 iovss.n2089 iovss.n2013 9.0005
R19 iovss.n2089 iovss.n2019 9.0005
R20 iovss.n2089 iovss.n2011 9.0005
R21 iovss.n2089 iovss.n2021 9.0005
R22 iovss.n2089 iovss.n2009 9.0005
R23 iovss.n2089 iovss.n2008 9.0005
R24 iovss.n2089 iovss.n2026 9.0005
R25 iovss.n2089 iovss.n2006 9.0005
R26 iovss.n2089 iovss.n2028 9.0005
R27 iovss.n2089 iovss.n2004 9.0005
R28 iovss.n2089 iovss.n2030 9.0005
R29 iovss.n2089 iovss.n2002 9.0005
R30 iovss.n2089 iovss.n2032 9.0005
R31 iovss.n2089 iovss.n2000 9.0005
R32 iovss.n2089 iovss.n2078 9.0005
R33 iovss.n2090 iovss.n2089 9.0005
R34 iovss.n2092 iovss.n1440 9.0005
R35 iovss.n2016 iovss.n1440 9.0005
R36 iovss.n2015 iovss.n1440 9.0005
R37 iovss.n2017 iovss.n1440 9.0005
R38 iovss.n2014 iovss.n1440 9.0005
R39 iovss.n2018 iovss.n1440 9.0005
R40 iovss.n2013 iovss.n1440 9.0005
R41 iovss.n2019 iovss.n1440 9.0005
R42 iovss.n2012 iovss.n1440 9.0005
R43 iovss.n2020 iovss.n1440 9.0005
R44 iovss.n2011 iovss.n1440 9.0005
R45 iovss.n2021 iovss.n1440 9.0005
R46 iovss.n2010 iovss.n1440 9.0005
R47 iovss.n2022 iovss.n1440 9.0005
R48 iovss.n2009 iovss.n1440 9.0005
R49 iovss.n2025 iovss.n1440 9.0005
R50 iovss.n2007 iovss.n1440 9.0005
R51 iovss.n2026 iovss.n1440 9.0005
R52 iovss.n2006 iovss.n1440 9.0005
R53 iovss.n2027 iovss.n1440 9.0005
R54 iovss.n2005 iovss.n1440 9.0005
R55 iovss.n2028 iovss.n1440 9.0005
R56 iovss.n2004 iovss.n1440 9.0005
R57 iovss.n2029 iovss.n1440 9.0005
R58 iovss.n2003 iovss.n1440 9.0005
R59 iovss.n2030 iovss.n1440 9.0005
R60 iovss.n2002 iovss.n1440 9.0005
R61 iovss.n2031 iovss.n1440 9.0005
R62 iovss.n2001 iovss.n1440 9.0005
R63 iovss.n2032 iovss.n1440 9.0005
R64 iovss.n2000 iovss.n1440 9.0005
R65 iovss.n2033 iovss.n1440 9.0005
R66 iovss.n2080 iovss.n1440 9.0005
R67 iovss.n2078 iovss.n1440 9.0005
R68 iovss.n2090 iovss.n1440 9.0005
R69 iovss.n2092 iovss.n1441 9.0005
R70 iovss.n2016 iovss.n1441 9.0005
R71 iovss.n2015 iovss.n1441 9.0005
R72 iovss.n2017 iovss.n1441 9.0005
R73 iovss.n2014 iovss.n1441 9.0005
R74 iovss.n2018 iovss.n1441 9.0005
R75 iovss.n2013 iovss.n1441 9.0005
R76 iovss.n2019 iovss.n1441 9.0005
R77 iovss.n2012 iovss.n1441 9.0005
R78 iovss.n2020 iovss.n1441 9.0005
R79 iovss.n2011 iovss.n1441 9.0005
R80 iovss.n2021 iovss.n1441 9.0005
R81 iovss.n2010 iovss.n1441 9.0005
R82 iovss.n2022 iovss.n1441 9.0005
R83 iovss.n2009 iovss.n1441 9.0005
R84 iovss.n2024 iovss.n1441 9.0005
R85 iovss.n2008 iovss.n1441 9.0005
R86 iovss.n2025 iovss.n1441 9.0005
R87 iovss.n2007 iovss.n1441 9.0005
R88 iovss.n2026 iovss.n1441 9.0005
R89 iovss.n2006 iovss.n1441 9.0005
R90 iovss.n2027 iovss.n1441 9.0005
R91 iovss.n2005 iovss.n1441 9.0005
R92 iovss.n2028 iovss.n1441 9.0005
R93 iovss.n2004 iovss.n1441 9.0005
R94 iovss.n2029 iovss.n1441 9.0005
R95 iovss.n2003 iovss.n1441 9.0005
R96 iovss.n2030 iovss.n1441 9.0005
R97 iovss.n2002 iovss.n1441 9.0005
R98 iovss.n2031 iovss.n1441 9.0005
R99 iovss.n2001 iovss.n1441 9.0005
R100 iovss.n2032 iovss.n1441 9.0005
R101 iovss.n2000 iovss.n1441 9.0005
R102 iovss.n2033 iovss.n1441 9.0005
R103 iovss.n2080 iovss.n1441 9.0005
R104 iovss.n2078 iovss.n1441 9.0005
R105 iovss.n2090 iovss.n1441 9.0005
R106 iovss.n2092 iovss.n1982 9.0005
R107 iovss.n2016 iovss.n1982 9.0005
R108 iovss.n2015 iovss.n1982 9.0005
R109 iovss.n2017 iovss.n1982 9.0005
R110 iovss.n2014 iovss.n1982 9.0005
R111 iovss.n2018 iovss.n1982 9.0005
R112 iovss.n2013 iovss.n1982 9.0005
R113 iovss.n2019 iovss.n1982 9.0005
R114 iovss.n2012 iovss.n1982 9.0005
R115 iovss.n2020 iovss.n1982 9.0005
R116 iovss.n2011 iovss.n1982 9.0005
R117 iovss.n2021 iovss.n1982 9.0005
R118 iovss.n2010 iovss.n1982 9.0005
R119 iovss.n2022 iovss.n1982 9.0005
R120 iovss.n2009 iovss.n1982 9.0005
R121 iovss.n2024 iovss.n1982 9.0005
R122 iovss.n2008 iovss.n1982 9.0005
R123 iovss.n2025 iovss.n1982 9.0005
R124 iovss.n2007 iovss.n1982 9.0005
R125 iovss.n2026 iovss.n1982 9.0005
R126 iovss.n2006 iovss.n1982 9.0005
R127 iovss.n2027 iovss.n1982 9.0005
R128 iovss.n2005 iovss.n1982 9.0005
R129 iovss.n2028 iovss.n1982 9.0005
R130 iovss.n2004 iovss.n1982 9.0005
R131 iovss.n2029 iovss.n1982 9.0005
R132 iovss.n2003 iovss.n1982 9.0005
R133 iovss.n2030 iovss.n1982 9.0005
R134 iovss.n2002 iovss.n1982 9.0005
R135 iovss.n2031 iovss.n1982 9.0005
R136 iovss.n2001 iovss.n1982 9.0005
R137 iovss.n2032 iovss.n1982 9.0005
R138 iovss.n2000 iovss.n1982 9.0005
R139 iovss.n2033 iovss.n1982 9.0005
R140 iovss.n2078 iovss.n1982 9.0005
R141 iovss.n2090 iovss.n1982 9.0005
R142 iovss.n2092 iovss.n2091 9.0005
R143 iovss.n2091 iovss.n2016 9.0005
R144 iovss.n2091 iovss.n2015 9.0005
R145 iovss.n2091 iovss.n2017 9.0005
R146 iovss.n2091 iovss.n2014 9.0005
R147 iovss.n2091 iovss.n2018 9.0005
R148 iovss.n2091 iovss.n2013 9.0005
R149 iovss.n2091 iovss.n2019 9.0005
R150 iovss.n2091 iovss.n2012 9.0005
R151 iovss.n2091 iovss.n2020 9.0005
R152 iovss.n2091 iovss.n2011 9.0005
R153 iovss.n2091 iovss.n2021 9.0005
R154 iovss.n2091 iovss.n2010 9.0005
R155 iovss.n2091 iovss.n2022 9.0005
R156 iovss.n2091 iovss.n2009 9.0005
R157 iovss.n2091 iovss.n2024 9.0005
R158 iovss.n2091 iovss.n2008 9.0005
R159 iovss.n2091 iovss.n2025 9.0005
R160 iovss.n2091 iovss.n2007 9.0005
R161 iovss.n2091 iovss.n2026 9.0005
R162 iovss.n2091 iovss.n2006 9.0005
R163 iovss.n2091 iovss.n2027 9.0005
R164 iovss.n2091 iovss.n2005 9.0005
R165 iovss.n2091 iovss.n2028 9.0005
R166 iovss.n2091 iovss.n2004 9.0005
R167 iovss.n2091 iovss.n2029 9.0005
R168 iovss.n2091 iovss.n2003 9.0005
R169 iovss.n2091 iovss.n2030 9.0005
R170 iovss.n2091 iovss.n2002 9.0005
R171 iovss.n2091 iovss.n2031 9.0005
R172 iovss.n2091 iovss.n2001 9.0005
R173 iovss.n2091 iovss.n2032 9.0005
R174 iovss.n2091 iovss.n2000 9.0005
R175 iovss.n2091 iovss.n2033 9.0005
R176 iovss.n2091 iovss.n2078 9.0005
R177 iovss.n2091 iovss.n1999 9.0005
R178 iovss.n2091 iovss.n2090 9.0005
R179 iovss.n1547 iovss.n1546 9.0005
R180 iovss.n1546 iovss.n1536 9.0005
R181 iovss.n1546 iovss.n1545 9.0005
R182 iovss.n1539 iovss.n1536 9.0005
R183 iovss.n1545 iovss.n1539 9.0005
R184 iovss.n1545 iovss.n1442 9.0005
R185 iovss.n1536 iovss.n1445 9.0005
R186 iovss.n1538 iovss.n1536 9.0005
R187 iovss.n1545 iovss.n1538 9.0005
R188 iovss.n1545 iovss.n1544 9.0005
R189 iovss.n1996 iovss.n1984 9.0005
R190 iovss.n1994 iovss.n1987 9.0005
R191 iovss.n1996 iovss.n1987 9.0005
R192 iovss.n1996 iovss.n1446 9.0005
R193 iovss.n1485 iovss.n1447 9.0005
R194 iovss.n1994 iovss.n1447 9.0005
R195 iovss.n1996 iovss.n1447 9.0005
R196 iovss.n1994 iovss.n1983 9.0005
R197 iovss.n1996 iovss.n1983 9.0005
R198 iovss.n1995 iovss.n1994 9.0005
R199 iovss.n1995 iovss.n1991 9.0005
R200 iovss.n1996 iovss.n1995 9.0005
R201 iovss.n1502 iovss.n1467 9.0005
R202 iovss.n1502 iovss.n1469 9.0005
R203 iovss.n1502 iovss.n1465 9.0005
R204 iovss.n2560 iovss.n1502 9.0005
R205 iovss.n2562 iovss.n1502 9.0005
R206 iovss.n2552 iovss.n1461 9.0005
R207 iovss.n2552 iovss.n1474 9.0005
R208 iovss.n2552 iovss.n1459 9.0005
R209 iovss.n2552 iovss.n1476 9.0005
R210 iovss.n2552 iovss.n1457 9.0005
R211 iovss.n2552 iovss.n1478 9.0005
R212 iovss.n2552 iovss.n1455 9.0005
R213 iovss.n2552 iovss.n1480 9.0005
R214 iovss.n2552 iovss.n1453 9.0005
R215 iovss.n2552 iovss.n1482 9.0005
R216 iovss.n2552 iovss.n1451 9.0005
R217 iovss.n2552 iovss.n1484 9.0005
R218 iovss.n2560 iovss.n2552 9.0005
R219 iovss.n2562 iovss.n2552 9.0005
R220 iovss.n1467 iovss.n1448 9.0005
R221 iovss.n1468 iovss.n1448 9.0005
R222 iovss.n1466 iovss.n1448 9.0005
R223 iovss.n1469 iovss.n1448 9.0005
R224 iovss.n1465 iovss.n1448 9.0005
R225 iovss.n1470 iovss.n1448 9.0005
R226 iovss.n1464 iovss.n1448 9.0005
R227 iovss.n1471 iovss.n1448 9.0005
R228 iovss.n1463 iovss.n1448 9.0005
R229 iovss.n1472 iovss.n1448 9.0005
R230 iovss.n1462 iovss.n1448 9.0005
R231 iovss.n1473 iovss.n1448 9.0005
R232 iovss.n1461 iovss.n1448 9.0005
R233 iovss.n1474 iovss.n1448 9.0005
R234 iovss.n1460 iovss.n1448 9.0005
R235 iovss.n1475 iovss.n1448 9.0005
R236 iovss.n1459 iovss.n1448 9.0005
R237 iovss.n1476 iovss.n1448 9.0005
R238 iovss.n1458 iovss.n1448 9.0005
R239 iovss.n1477 iovss.n1448 9.0005
R240 iovss.n1457 iovss.n1448 9.0005
R241 iovss.n1478 iovss.n1448 9.0005
R242 iovss.n1456 iovss.n1448 9.0005
R243 iovss.n1479 iovss.n1448 9.0005
R244 iovss.n1455 iovss.n1448 9.0005
R245 iovss.n1480 iovss.n1448 9.0005
R246 iovss.n1454 iovss.n1448 9.0005
R247 iovss.n1481 iovss.n1448 9.0005
R248 iovss.n1453 iovss.n1448 9.0005
R249 iovss.n1482 iovss.n1448 9.0005
R250 iovss.n1452 iovss.n1448 9.0005
R251 iovss.n1483 iovss.n1448 9.0005
R252 iovss.n1451 iovss.n1448 9.0005
R253 iovss.n1484 iovss.n1448 9.0005
R254 iovss.n2562 iovss.n1448 9.0005
R255 iovss.n2563 iovss.n1467 9.0005
R256 iovss.n2563 iovss.n1468 9.0005
R257 iovss.n2563 iovss.n1466 9.0005
R258 iovss.n2563 iovss.n1469 9.0005
R259 iovss.n2563 iovss.n1465 9.0005
R260 iovss.n2563 iovss.n1470 9.0005
R261 iovss.n2563 iovss.n1464 9.0005
R262 iovss.n2563 iovss.n1471 9.0005
R263 iovss.n2563 iovss.n1463 9.0005
R264 iovss.n2563 iovss.n1472 9.0005
R265 iovss.n2563 iovss.n1462 9.0005
R266 iovss.n2563 iovss.n1473 9.0005
R267 iovss.n2563 iovss.n1461 9.0005
R268 iovss.n2563 iovss.n1474 9.0005
R269 iovss.n2563 iovss.n1460 9.0005
R270 iovss.n2563 iovss.n1475 9.0005
R271 iovss.n2563 iovss.n1459 9.0005
R272 iovss.n2563 iovss.n1476 9.0005
R273 iovss.n2563 iovss.n1458 9.0005
R274 iovss.n2563 iovss.n1477 9.0005
R275 iovss.n2563 iovss.n1457 9.0005
R276 iovss.n2563 iovss.n1478 9.0005
R277 iovss.n2563 iovss.n1456 9.0005
R278 iovss.n2563 iovss.n1479 9.0005
R279 iovss.n2563 iovss.n1455 9.0005
R280 iovss.n2563 iovss.n1480 9.0005
R281 iovss.n2563 iovss.n1454 9.0005
R282 iovss.n2563 iovss.n1481 9.0005
R283 iovss.n2563 iovss.n1453 9.0005
R284 iovss.n2563 iovss.n1482 9.0005
R285 iovss.n2563 iovss.n1452 9.0005
R286 iovss.n2563 iovss.n1483 9.0005
R287 iovss.n2563 iovss.n1451 9.0005
R288 iovss.n2563 iovss.n1484 9.0005
R289 iovss.n2563 iovss.n2562 9.0005
R290 iovss.n1486 iovss.n1467 9.0005
R291 iovss.n1486 iovss.n1468 9.0005
R292 iovss.n1486 iovss.n1466 9.0005
R293 iovss.n1486 iovss.n1469 9.0005
R294 iovss.n1486 iovss.n1465 9.0005
R295 iovss.n1486 iovss.n1470 9.0005
R296 iovss.n1486 iovss.n1464 9.0005
R297 iovss.n1486 iovss.n1471 9.0005
R298 iovss.n1486 iovss.n1463 9.0005
R299 iovss.n1486 iovss.n1472 9.0005
R300 iovss.n1486 iovss.n1462 9.0005
R301 iovss.n1486 iovss.n1473 9.0005
R302 iovss.n1486 iovss.n1461 9.0005
R303 iovss.n1486 iovss.n1474 9.0005
R304 iovss.n1486 iovss.n1460 9.0005
R305 iovss.n1486 iovss.n1475 9.0005
R306 iovss.n1486 iovss.n1459 9.0005
R307 iovss.n1486 iovss.n1476 9.0005
R308 iovss.n1486 iovss.n1458 9.0005
R309 iovss.n1486 iovss.n1477 9.0005
R310 iovss.n1486 iovss.n1457 9.0005
R311 iovss.n1486 iovss.n1478 9.0005
R312 iovss.n1486 iovss.n1456 9.0005
R313 iovss.n1486 iovss.n1479 9.0005
R314 iovss.n1486 iovss.n1455 9.0005
R315 iovss.n1486 iovss.n1480 9.0005
R316 iovss.n1486 iovss.n1454 9.0005
R317 iovss.n1486 iovss.n1481 9.0005
R318 iovss.n1486 iovss.n1453 9.0005
R319 iovss.n1486 iovss.n1482 9.0005
R320 iovss.n1486 iovss.n1452 9.0005
R321 iovss.n1486 iovss.n1483 9.0005
R322 iovss.n1486 iovss.n1451 9.0005
R323 iovss.n1486 iovss.n1484 9.0005
R324 iovss.n2560 iovss.n1486 9.0005
R325 iovss.n2562 iovss.n1486 9.0005
R326 iovss.n2561 iovss.n1467 9.0005
R327 iovss.n2561 iovss.n1468 9.0005
R328 iovss.n2561 iovss.n1466 9.0005
R329 iovss.n2561 iovss.n1469 9.0005
R330 iovss.n2561 iovss.n1465 9.0005
R331 iovss.n2561 iovss.n1470 9.0005
R332 iovss.n2561 iovss.n1464 9.0005
R333 iovss.n2561 iovss.n1471 9.0005
R334 iovss.n2561 iovss.n1463 9.0005
R335 iovss.n2561 iovss.n1472 9.0005
R336 iovss.n2561 iovss.n1462 9.0005
R337 iovss.n2561 iovss.n1473 9.0005
R338 iovss.n2561 iovss.n1461 9.0005
R339 iovss.n2561 iovss.n1474 9.0005
R340 iovss.n2561 iovss.n1460 9.0005
R341 iovss.n2561 iovss.n1475 9.0005
R342 iovss.n2561 iovss.n1459 9.0005
R343 iovss.n2561 iovss.n1476 9.0005
R344 iovss.n2561 iovss.n1458 9.0005
R345 iovss.n2561 iovss.n1477 9.0005
R346 iovss.n2561 iovss.n1457 9.0005
R347 iovss.n2561 iovss.n1478 9.0005
R348 iovss.n2561 iovss.n1456 9.0005
R349 iovss.n2561 iovss.n1479 9.0005
R350 iovss.n2561 iovss.n1455 9.0005
R351 iovss.n2561 iovss.n1480 9.0005
R352 iovss.n2561 iovss.n1454 9.0005
R353 iovss.n2561 iovss.n1481 9.0005
R354 iovss.n2561 iovss.n1453 9.0005
R355 iovss.n2561 iovss.n1482 9.0005
R356 iovss.n2561 iovss.n1452 9.0005
R357 iovss.n2561 iovss.n1483 9.0005
R358 iovss.n2561 iovss.n1451 9.0005
R359 iovss.n2561 iovss.n1484 9.0005
R360 iovss.n2561 iovss.n2560 9.0005
R361 iovss.n2561 iovss.n2558 9.0005
R362 iovss.n2562 iovss.n2561 9.0005
R363 iovss.n1790 iovss.n303 9.0005
R364 iovss.n2292 iovss.n1732 9.0005
R365 iovss.n1804 iovss.n1732 9.0005
R366 iovss.n1798 iovss.n1732 9.0005
R367 iovss.n1809 iovss.n1732 9.0005
R368 iovss.n1796 iovss.n1732 9.0005
R369 iovss.n1814 iovss.n1732 9.0005
R370 iovss.n1794 iovss.n1732 9.0005
R371 iovss.n1819 iovss.n1732 9.0005
R372 iovss.n1792 iovss.n1732 9.0005
R373 iovss.n1824 iovss.n1732 9.0005
R374 iovss.n1788 iovss.n1732 9.0005
R375 iovss.n1832 iovss.n1732 9.0005
R376 iovss.n1786 iovss.n1732 9.0005
R377 iovss.n1837 iovss.n1732 9.0005
R378 iovss.n1784 iovss.n1732 9.0005
R379 iovss.n1841 iovss.n1732 9.0005
R380 iovss.n2292 iovss.n1730 9.0005
R381 iovss.n1801 iovss.n1730 9.0005
R382 iovss.n1799 iovss.n1730 9.0005
R383 iovss.n1804 iovss.n1730 9.0005
R384 iovss.n1798 iovss.n1730 9.0005
R385 iovss.n1807 iovss.n1730 9.0005
R386 iovss.n1797 iovss.n1730 9.0005
R387 iovss.n1809 iovss.n1730 9.0005
R388 iovss.n1796 iovss.n1730 9.0005
R389 iovss.n1812 iovss.n1730 9.0005
R390 iovss.n1795 iovss.n1730 9.0005
R391 iovss.n1814 iovss.n1730 9.0005
R392 iovss.n1794 iovss.n1730 9.0005
R393 iovss.n1817 iovss.n1730 9.0005
R394 iovss.n1793 iovss.n1730 9.0005
R395 iovss.n1819 iovss.n1730 9.0005
R396 iovss.n1792 iovss.n1730 9.0005
R397 iovss.n1822 iovss.n1730 9.0005
R398 iovss.n1791 iovss.n1730 9.0005
R399 iovss.n1824 iovss.n1730 9.0005
R400 iovss.n1790 iovss.n1730 9.0005
R401 iovss.n1827 iovss.n1730 9.0005
R402 iovss.n1789 iovss.n1730 9.0005
R403 iovss.n1830 iovss.n1730 9.0005
R404 iovss.n1788 iovss.n1730 9.0005
R405 iovss.n1832 iovss.n1730 9.0005
R406 iovss.n1787 iovss.n1730 9.0005
R407 iovss.n1835 iovss.n1730 9.0005
R408 iovss.n1786 iovss.n1730 9.0005
R409 iovss.n1837 iovss.n1730 9.0005
R410 iovss.n1785 iovss.n1730 9.0005
R411 iovss.n1840 iovss.n1730 9.0005
R412 iovss.n1784 iovss.n1730 9.0005
R413 iovss.n1841 iovss.n1730 9.0005
R414 iovss.n1870 iovss.n1730 9.0005
R415 iovss.n2290 iovss.n1730 9.0005
R416 iovss.n2292 iovss.n1733 9.0005
R417 iovss.n1801 iovss.n1733 9.0005
R418 iovss.n1799 iovss.n1733 9.0005
R419 iovss.n1804 iovss.n1733 9.0005
R420 iovss.n1798 iovss.n1733 9.0005
R421 iovss.n1807 iovss.n1733 9.0005
R422 iovss.n1797 iovss.n1733 9.0005
R423 iovss.n1809 iovss.n1733 9.0005
R424 iovss.n1796 iovss.n1733 9.0005
R425 iovss.n1812 iovss.n1733 9.0005
R426 iovss.n1795 iovss.n1733 9.0005
R427 iovss.n1814 iovss.n1733 9.0005
R428 iovss.n1794 iovss.n1733 9.0005
R429 iovss.n1817 iovss.n1733 9.0005
R430 iovss.n1793 iovss.n1733 9.0005
R431 iovss.n1819 iovss.n1733 9.0005
R432 iovss.n1792 iovss.n1733 9.0005
R433 iovss.n1822 iovss.n1733 9.0005
R434 iovss.n1791 iovss.n1733 9.0005
R435 iovss.n1824 iovss.n1733 9.0005
R436 iovss.n1790 iovss.n1733 9.0005
R437 iovss.n1827 iovss.n1733 9.0005
R438 iovss.n1789 iovss.n1733 9.0005
R439 iovss.n1830 iovss.n1733 9.0005
R440 iovss.n1788 iovss.n1733 9.0005
R441 iovss.n1832 iovss.n1733 9.0005
R442 iovss.n1787 iovss.n1733 9.0005
R443 iovss.n1835 iovss.n1733 9.0005
R444 iovss.n1786 iovss.n1733 9.0005
R445 iovss.n1837 iovss.n1733 9.0005
R446 iovss.n1785 iovss.n1733 9.0005
R447 iovss.n1840 iovss.n1733 9.0005
R448 iovss.n1784 iovss.n1733 9.0005
R449 iovss.n1841 iovss.n1733 9.0005
R450 iovss.n1870 iovss.n1733 9.0005
R451 iovss.n2290 iovss.n1733 9.0005
R452 iovss.n2292 iovss.n1729 9.0005
R453 iovss.n1801 iovss.n1729 9.0005
R454 iovss.n1799 iovss.n1729 9.0005
R455 iovss.n1804 iovss.n1729 9.0005
R456 iovss.n1798 iovss.n1729 9.0005
R457 iovss.n1807 iovss.n1729 9.0005
R458 iovss.n1797 iovss.n1729 9.0005
R459 iovss.n1809 iovss.n1729 9.0005
R460 iovss.n1796 iovss.n1729 9.0005
R461 iovss.n1812 iovss.n1729 9.0005
R462 iovss.n1795 iovss.n1729 9.0005
R463 iovss.n1814 iovss.n1729 9.0005
R464 iovss.n1794 iovss.n1729 9.0005
R465 iovss.n1817 iovss.n1729 9.0005
R466 iovss.n1793 iovss.n1729 9.0005
R467 iovss.n1819 iovss.n1729 9.0005
R468 iovss.n1792 iovss.n1729 9.0005
R469 iovss.n1822 iovss.n1729 9.0005
R470 iovss.n1791 iovss.n1729 9.0005
R471 iovss.n1824 iovss.n1729 9.0005
R472 iovss.n1790 iovss.n1729 9.0005
R473 iovss.n1827 iovss.n1729 9.0005
R474 iovss.n1789 iovss.n1729 9.0005
R475 iovss.n1830 iovss.n1729 9.0005
R476 iovss.n1788 iovss.n1729 9.0005
R477 iovss.n1832 iovss.n1729 9.0005
R478 iovss.n1787 iovss.n1729 9.0005
R479 iovss.n1835 iovss.n1729 9.0005
R480 iovss.n1786 iovss.n1729 9.0005
R481 iovss.n1837 iovss.n1729 9.0005
R482 iovss.n1785 iovss.n1729 9.0005
R483 iovss.n1840 iovss.n1729 9.0005
R484 iovss.n1784 iovss.n1729 9.0005
R485 iovss.n1841 iovss.n1729 9.0005
R486 iovss.n1870 iovss.n1729 9.0005
R487 iovss.n2290 iovss.n1729 9.0005
R488 iovss.n2292 iovss.n1734 9.0005
R489 iovss.n1801 iovss.n1734 9.0005
R490 iovss.n1799 iovss.n1734 9.0005
R491 iovss.n1804 iovss.n1734 9.0005
R492 iovss.n1798 iovss.n1734 9.0005
R493 iovss.n1807 iovss.n1734 9.0005
R494 iovss.n1797 iovss.n1734 9.0005
R495 iovss.n1809 iovss.n1734 9.0005
R496 iovss.n1796 iovss.n1734 9.0005
R497 iovss.n1812 iovss.n1734 9.0005
R498 iovss.n1795 iovss.n1734 9.0005
R499 iovss.n1814 iovss.n1734 9.0005
R500 iovss.n1794 iovss.n1734 9.0005
R501 iovss.n1817 iovss.n1734 9.0005
R502 iovss.n1793 iovss.n1734 9.0005
R503 iovss.n1819 iovss.n1734 9.0005
R504 iovss.n1792 iovss.n1734 9.0005
R505 iovss.n1822 iovss.n1734 9.0005
R506 iovss.n1791 iovss.n1734 9.0005
R507 iovss.n1824 iovss.n1734 9.0005
R508 iovss.n1790 iovss.n1734 9.0005
R509 iovss.n1827 iovss.n1734 9.0005
R510 iovss.n1789 iovss.n1734 9.0005
R511 iovss.n1830 iovss.n1734 9.0005
R512 iovss.n1788 iovss.n1734 9.0005
R513 iovss.n1832 iovss.n1734 9.0005
R514 iovss.n1787 iovss.n1734 9.0005
R515 iovss.n1835 iovss.n1734 9.0005
R516 iovss.n1786 iovss.n1734 9.0005
R517 iovss.n1837 iovss.n1734 9.0005
R518 iovss.n1785 iovss.n1734 9.0005
R519 iovss.n1840 iovss.n1734 9.0005
R520 iovss.n1784 iovss.n1734 9.0005
R521 iovss.n1841 iovss.n1734 9.0005
R522 iovss.n1870 iovss.n1734 9.0005
R523 iovss.n2290 iovss.n1734 9.0005
R524 iovss.n2292 iovss.n1728 9.0005
R525 iovss.n1801 iovss.n1728 9.0005
R526 iovss.n1799 iovss.n1728 9.0005
R527 iovss.n1804 iovss.n1728 9.0005
R528 iovss.n1798 iovss.n1728 9.0005
R529 iovss.n1807 iovss.n1728 9.0005
R530 iovss.n1797 iovss.n1728 9.0005
R531 iovss.n1809 iovss.n1728 9.0005
R532 iovss.n1796 iovss.n1728 9.0005
R533 iovss.n1812 iovss.n1728 9.0005
R534 iovss.n1795 iovss.n1728 9.0005
R535 iovss.n1814 iovss.n1728 9.0005
R536 iovss.n1794 iovss.n1728 9.0005
R537 iovss.n1817 iovss.n1728 9.0005
R538 iovss.n1793 iovss.n1728 9.0005
R539 iovss.n1819 iovss.n1728 9.0005
R540 iovss.n1792 iovss.n1728 9.0005
R541 iovss.n1822 iovss.n1728 9.0005
R542 iovss.n1791 iovss.n1728 9.0005
R543 iovss.n1824 iovss.n1728 9.0005
R544 iovss.n1790 iovss.n1728 9.0005
R545 iovss.n1827 iovss.n1728 9.0005
R546 iovss.n1789 iovss.n1728 9.0005
R547 iovss.n1830 iovss.n1728 9.0005
R548 iovss.n1788 iovss.n1728 9.0005
R549 iovss.n1832 iovss.n1728 9.0005
R550 iovss.n1787 iovss.n1728 9.0005
R551 iovss.n1835 iovss.n1728 9.0005
R552 iovss.n1786 iovss.n1728 9.0005
R553 iovss.n1837 iovss.n1728 9.0005
R554 iovss.n1785 iovss.n1728 9.0005
R555 iovss.n1840 iovss.n1728 9.0005
R556 iovss.n1784 iovss.n1728 9.0005
R557 iovss.n1841 iovss.n1728 9.0005
R558 iovss.n1870 iovss.n1728 9.0005
R559 iovss.n2290 iovss.n1728 9.0005
R560 iovss.n2292 iovss.n1735 9.0005
R561 iovss.n1801 iovss.n1735 9.0005
R562 iovss.n1799 iovss.n1735 9.0005
R563 iovss.n1804 iovss.n1735 9.0005
R564 iovss.n1798 iovss.n1735 9.0005
R565 iovss.n1807 iovss.n1735 9.0005
R566 iovss.n1797 iovss.n1735 9.0005
R567 iovss.n1809 iovss.n1735 9.0005
R568 iovss.n1796 iovss.n1735 9.0005
R569 iovss.n1812 iovss.n1735 9.0005
R570 iovss.n1795 iovss.n1735 9.0005
R571 iovss.n1814 iovss.n1735 9.0005
R572 iovss.n1794 iovss.n1735 9.0005
R573 iovss.n1817 iovss.n1735 9.0005
R574 iovss.n1793 iovss.n1735 9.0005
R575 iovss.n1819 iovss.n1735 9.0005
R576 iovss.n1792 iovss.n1735 9.0005
R577 iovss.n1822 iovss.n1735 9.0005
R578 iovss.n1791 iovss.n1735 9.0005
R579 iovss.n1824 iovss.n1735 9.0005
R580 iovss.n1790 iovss.n1735 9.0005
R581 iovss.n1827 iovss.n1735 9.0005
R582 iovss.n1789 iovss.n1735 9.0005
R583 iovss.n1830 iovss.n1735 9.0005
R584 iovss.n1788 iovss.n1735 9.0005
R585 iovss.n1832 iovss.n1735 9.0005
R586 iovss.n1787 iovss.n1735 9.0005
R587 iovss.n1835 iovss.n1735 9.0005
R588 iovss.n1786 iovss.n1735 9.0005
R589 iovss.n1837 iovss.n1735 9.0005
R590 iovss.n1785 iovss.n1735 9.0005
R591 iovss.n1840 iovss.n1735 9.0005
R592 iovss.n1784 iovss.n1735 9.0005
R593 iovss.n1841 iovss.n1735 9.0005
R594 iovss.n1870 iovss.n1735 9.0005
R595 iovss.n2290 iovss.n1735 9.0005
R596 iovss.n2292 iovss.n1727 9.0005
R597 iovss.n1801 iovss.n1727 9.0005
R598 iovss.n1799 iovss.n1727 9.0005
R599 iovss.n1804 iovss.n1727 9.0005
R600 iovss.n1798 iovss.n1727 9.0005
R601 iovss.n1807 iovss.n1727 9.0005
R602 iovss.n1797 iovss.n1727 9.0005
R603 iovss.n1809 iovss.n1727 9.0005
R604 iovss.n1796 iovss.n1727 9.0005
R605 iovss.n1812 iovss.n1727 9.0005
R606 iovss.n1795 iovss.n1727 9.0005
R607 iovss.n1814 iovss.n1727 9.0005
R608 iovss.n1794 iovss.n1727 9.0005
R609 iovss.n1817 iovss.n1727 9.0005
R610 iovss.n1793 iovss.n1727 9.0005
R611 iovss.n1819 iovss.n1727 9.0005
R612 iovss.n1792 iovss.n1727 9.0005
R613 iovss.n1822 iovss.n1727 9.0005
R614 iovss.n1791 iovss.n1727 9.0005
R615 iovss.n1824 iovss.n1727 9.0005
R616 iovss.n1790 iovss.n1727 9.0005
R617 iovss.n1827 iovss.n1727 9.0005
R618 iovss.n1789 iovss.n1727 9.0005
R619 iovss.n1830 iovss.n1727 9.0005
R620 iovss.n1788 iovss.n1727 9.0005
R621 iovss.n1832 iovss.n1727 9.0005
R622 iovss.n1787 iovss.n1727 9.0005
R623 iovss.n1835 iovss.n1727 9.0005
R624 iovss.n1786 iovss.n1727 9.0005
R625 iovss.n1837 iovss.n1727 9.0005
R626 iovss.n1785 iovss.n1727 9.0005
R627 iovss.n1840 iovss.n1727 9.0005
R628 iovss.n1784 iovss.n1727 9.0005
R629 iovss.n1841 iovss.n1727 9.0005
R630 iovss.n1870 iovss.n1727 9.0005
R631 iovss.n2290 iovss.n1727 9.0005
R632 iovss.n2292 iovss.n1736 9.0005
R633 iovss.n1801 iovss.n1736 9.0005
R634 iovss.n1799 iovss.n1736 9.0005
R635 iovss.n1804 iovss.n1736 9.0005
R636 iovss.n1798 iovss.n1736 9.0005
R637 iovss.n1807 iovss.n1736 9.0005
R638 iovss.n1797 iovss.n1736 9.0005
R639 iovss.n1809 iovss.n1736 9.0005
R640 iovss.n1796 iovss.n1736 9.0005
R641 iovss.n1812 iovss.n1736 9.0005
R642 iovss.n1795 iovss.n1736 9.0005
R643 iovss.n1814 iovss.n1736 9.0005
R644 iovss.n1794 iovss.n1736 9.0005
R645 iovss.n1817 iovss.n1736 9.0005
R646 iovss.n1793 iovss.n1736 9.0005
R647 iovss.n1819 iovss.n1736 9.0005
R648 iovss.n1792 iovss.n1736 9.0005
R649 iovss.n1822 iovss.n1736 9.0005
R650 iovss.n1791 iovss.n1736 9.0005
R651 iovss.n1824 iovss.n1736 9.0005
R652 iovss.n1790 iovss.n1736 9.0005
R653 iovss.n1827 iovss.n1736 9.0005
R654 iovss.n1789 iovss.n1736 9.0005
R655 iovss.n1830 iovss.n1736 9.0005
R656 iovss.n1788 iovss.n1736 9.0005
R657 iovss.n1832 iovss.n1736 9.0005
R658 iovss.n1787 iovss.n1736 9.0005
R659 iovss.n1835 iovss.n1736 9.0005
R660 iovss.n1786 iovss.n1736 9.0005
R661 iovss.n1837 iovss.n1736 9.0005
R662 iovss.n1785 iovss.n1736 9.0005
R663 iovss.n1840 iovss.n1736 9.0005
R664 iovss.n1784 iovss.n1736 9.0005
R665 iovss.n1841 iovss.n1736 9.0005
R666 iovss.n1870 iovss.n1736 9.0005
R667 iovss.n2290 iovss.n1736 9.0005
R668 iovss.n2292 iovss.n1726 9.0005
R669 iovss.n1801 iovss.n1726 9.0005
R670 iovss.n1799 iovss.n1726 9.0005
R671 iovss.n1804 iovss.n1726 9.0005
R672 iovss.n1798 iovss.n1726 9.0005
R673 iovss.n1807 iovss.n1726 9.0005
R674 iovss.n1797 iovss.n1726 9.0005
R675 iovss.n1809 iovss.n1726 9.0005
R676 iovss.n1796 iovss.n1726 9.0005
R677 iovss.n1812 iovss.n1726 9.0005
R678 iovss.n1795 iovss.n1726 9.0005
R679 iovss.n1814 iovss.n1726 9.0005
R680 iovss.n1794 iovss.n1726 9.0005
R681 iovss.n1817 iovss.n1726 9.0005
R682 iovss.n1793 iovss.n1726 9.0005
R683 iovss.n1819 iovss.n1726 9.0005
R684 iovss.n1792 iovss.n1726 9.0005
R685 iovss.n1822 iovss.n1726 9.0005
R686 iovss.n1791 iovss.n1726 9.0005
R687 iovss.n1824 iovss.n1726 9.0005
R688 iovss.n1790 iovss.n1726 9.0005
R689 iovss.n1827 iovss.n1726 9.0005
R690 iovss.n1789 iovss.n1726 9.0005
R691 iovss.n1830 iovss.n1726 9.0005
R692 iovss.n1788 iovss.n1726 9.0005
R693 iovss.n1832 iovss.n1726 9.0005
R694 iovss.n1787 iovss.n1726 9.0005
R695 iovss.n1835 iovss.n1726 9.0005
R696 iovss.n1786 iovss.n1726 9.0005
R697 iovss.n1837 iovss.n1726 9.0005
R698 iovss.n1785 iovss.n1726 9.0005
R699 iovss.n1840 iovss.n1726 9.0005
R700 iovss.n1784 iovss.n1726 9.0005
R701 iovss.n1841 iovss.n1726 9.0005
R702 iovss.n1870 iovss.n1726 9.0005
R703 iovss.n2290 iovss.n1726 9.0005
R704 iovss.n2292 iovss.n1737 9.0005
R705 iovss.n1801 iovss.n1737 9.0005
R706 iovss.n1799 iovss.n1737 9.0005
R707 iovss.n1804 iovss.n1737 9.0005
R708 iovss.n1798 iovss.n1737 9.0005
R709 iovss.n1807 iovss.n1737 9.0005
R710 iovss.n1797 iovss.n1737 9.0005
R711 iovss.n1809 iovss.n1737 9.0005
R712 iovss.n1796 iovss.n1737 9.0005
R713 iovss.n1812 iovss.n1737 9.0005
R714 iovss.n1795 iovss.n1737 9.0005
R715 iovss.n1814 iovss.n1737 9.0005
R716 iovss.n1794 iovss.n1737 9.0005
R717 iovss.n1817 iovss.n1737 9.0005
R718 iovss.n1793 iovss.n1737 9.0005
R719 iovss.n1819 iovss.n1737 9.0005
R720 iovss.n1792 iovss.n1737 9.0005
R721 iovss.n1822 iovss.n1737 9.0005
R722 iovss.n1791 iovss.n1737 9.0005
R723 iovss.n1824 iovss.n1737 9.0005
R724 iovss.n1790 iovss.n1737 9.0005
R725 iovss.n1827 iovss.n1737 9.0005
R726 iovss.n1789 iovss.n1737 9.0005
R727 iovss.n1830 iovss.n1737 9.0005
R728 iovss.n1788 iovss.n1737 9.0005
R729 iovss.n1832 iovss.n1737 9.0005
R730 iovss.n1787 iovss.n1737 9.0005
R731 iovss.n1835 iovss.n1737 9.0005
R732 iovss.n1786 iovss.n1737 9.0005
R733 iovss.n1837 iovss.n1737 9.0005
R734 iovss.n1785 iovss.n1737 9.0005
R735 iovss.n1840 iovss.n1737 9.0005
R736 iovss.n1784 iovss.n1737 9.0005
R737 iovss.n1841 iovss.n1737 9.0005
R738 iovss.n1870 iovss.n1737 9.0005
R739 iovss.n2290 iovss.n1737 9.0005
R740 iovss.n2292 iovss.n1725 9.0005
R741 iovss.n1801 iovss.n1725 9.0005
R742 iovss.n1799 iovss.n1725 9.0005
R743 iovss.n1804 iovss.n1725 9.0005
R744 iovss.n1798 iovss.n1725 9.0005
R745 iovss.n1807 iovss.n1725 9.0005
R746 iovss.n1797 iovss.n1725 9.0005
R747 iovss.n1809 iovss.n1725 9.0005
R748 iovss.n1796 iovss.n1725 9.0005
R749 iovss.n1812 iovss.n1725 9.0005
R750 iovss.n1795 iovss.n1725 9.0005
R751 iovss.n1814 iovss.n1725 9.0005
R752 iovss.n1794 iovss.n1725 9.0005
R753 iovss.n1817 iovss.n1725 9.0005
R754 iovss.n1793 iovss.n1725 9.0005
R755 iovss.n1819 iovss.n1725 9.0005
R756 iovss.n1792 iovss.n1725 9.0005
R757 iovss.n1822 iovss.n1725 9.0005
R758 iovss.n1791 iovss.n1725 9.0005
R759 iovss.n1824 iovss.n1725 9.0005
R760 iovss.n1790 iovss.n1725 9.0005
R761 iovss.n1827 iovss.n1725 9.0005
R762 iovss.n1789 iovss.n1725 9.0005
R763 iovss.n1830 iovss.n1725 9.0005
R764 iovss.n1788 iovss.n1725 9.0005
R765 iovss.n1832 iovss.n1725 9.0005
R766 iovss.n1787 iovss.n1725 9.0005
R767 iovss.n1835 iovss.n1725 9.0005
R768 iovss.n1786 iovss.n1725 9.0005
R769 iovss.n1837 iovss.n1725 9.0005
R770 iovss.n1785 iovss.n1725 9.0005
R771 iovss.n1840 iovss.n1725 9.0005
R772 iovss.n1784 iovss.n1725 9.0005
R773 iovss.n1841 iovss.n1725 9.0005
R774 iovss.n1870 iovss.n1725 9.0005
R775 iovss.n2290 iovss.n1725 9.0005
R776 iovss.n2292 iovss.n1738 9.0005
R777 iovss.n1801 iovss.n1738 9.0005
R778 iovss.n1799 iovss.n1738 9.0005
R779 iovss.n1804 iovss.n1738 9.0005
R780 iovss.n1798 iovss.n1738 9.0005
R781 iovss.n1807 iovss.n1738 9.0005
R782 iovss.n1797 iovss.n1738 9.0005
R783 iovss.n1809 iovss.n1738 9.0005
R784 iovss.n1796 iovss.n1738 9.0005
R785 iovss.n1812 iovss.n1738 9.0005
R786 iovss.n1795 iovss.n1738 9.0005
R787 iovss.n1814 iovss.n1738 9.0005
R788 iovss.n1794 iovss.n1738 9.0005
R789 iovss.n1817 iovss.n1738 9.0005
R790 iovss.n1793 iovss.n1738 9.0005
R791 iovss.n1819 iovss.n1738 9.0005
R792 iovss.n1792 iovss.n1738 9.0005
R793 iovss.n1822 iovss.n1738 9.0005
R794 iovss.n1791 iovss.n1738 9.0005
R795 iovss.n1824 iovss.n1738 9.0005
R796 iovss.n1790 iovss.n1738 9.0005
R797 iovss.n1827 iovss.n1738 9.0005
R798 iovss.n1789 iovss.n1738 9.0005
R799 iovss.n1830 iovss.n1738 9.0005
R800 iovss.n1788 iovss.n1738 9.0005
R801 iovss.n1832 iovss.n1738 9.0005
R802 iovss.n1787 iovss.n1738 9.0005
R803 iovss.n1835 iovss.n1738 9.0005
R804 iovss.n1786 iovss.n1738 9.0005
R805 iovss.n1837 iovss.n1738 9.0005
R806 iovss.n1785 iovss.n1738 9.0005
R807 iovss.n1840 iovss.n1738 9.0005
R808 iovss.n1784 iovss.n1738 9.0005
R809 iovss.n1841 iovss.n1738 9.0005
R810 iovss.n1870 iovss.n1738 9.0005
R811 iovss.n2290 iovss.n1738 9.0005
R812 iovss.n2292 iovss.n1724 9.0005
R813 iovss.n1801 iovss.n1724 9.0005
R814 iovss.n1799 iovss.n1724 9.0005
R815 iovss.n1804 iovss.n1724 9.0005
R816 iovss.n1798 iovss.n1724 9.0005
R817 iovss.n1807 iovss.n1724 9.0005
R818 iovss.n1797 iovss.n1724 9.0005
R819 iovss.n1809 iovss.n1724 9.0005
R820 iovss.n1796 iovss.n1724 9.0005
R821 iovss.n1812 iovss.n1724 9.0005
R822 iovss.n1795 iovss.n1724 9.0005
R823 iovss.n1814 iovss.n1724 9.0005
R824 iovss.n1794 iovss.n1724 9.0005
R825 iovss.n1817 iovss.n1724 9.0005
R826 iovss.n1793 iovss.n1724 9.0005
R827 iovss.n1819 iovss.n1724 9.0005
R828 iovss.n1792 iovss.n1724 9.0005
R829 iovss.n1822 iovss.n1724 9.0005
R830 iovss.n1791 iovss.n1724 9.0005
R831 iovss.n1824 iovss.n1724 9.0005
R832 iovss.n1790 iovss.n1724 9.0005
R833 iovss.n1827 iovss.n1724 9.0005
R834 iovss.n1789 iovss.n1724 9.0005
R835 iovss.n1830 iovss.n1724 9.0005
R836 iovss.n1788 iovss.n1724 9.0005
R837 iovss.n1832 iovss.n1724 9.0005
R838 iovss.n1787 iovss.n1724 9.0005
R839 iovss.n1835 iovss.n1724 9.0005
R840 iovss.n1786 iovss.n1724 9.0005
R841 iovss.n1837 iovss.n1724 9.0005
R842 iovss.n1785 iovss.n1724 9.0005
R843 iovss.n1840 iovss.n1724 9.0005
R844 iovss.n1784 iovss.n1724 9.0005
R845 iovss.n1841 iovss.n1724 9.0005
R846 iovss.n1870 iovss.n1724 9.0005
R847 iovss.n2290 iovss.n1724 9.0005
R848 iovss.n2292 iovss.n1739 9.0005
R849 iovss.n1801 iovss.n1739 9.0005
R850 iovss.n1799 iovss.n1739 9.0005
R851 iovss.n1804 iovss.n1739 9.0005
R852 iovss.n1798 iovss.n1739 9.0005
R853 iovss.n1807 iovss.n1739 9.0005
R854 iovss.n1797 iovss.n1739 9.0005
R855 iovss.n1809 iovss.n1739 9.0005
R856 iovss.n1796 iovss.n1739 9.0005
R857 iovss.n1812 iovss.n1739 9.0005
R858 iovss.n1795 iovss.n1739 9.0005
R859 iovss.n1814 iovss.n1739 9.0005
R860 iovss.n1794 iovss.n1739 9.0005
R861 iovss.n1817 iovss.n1739 9.0005
R862 iovss.n1793 iovss.n1739 9.0005
R863 iovss.n1819 iovss.n1739 9.0005
R864 iovss.n1792 iovss.n1739 9.0005
R865 iovss.n1822 iovss.n1739 9.0005
R866 iovss.n1791 iovss.n1739 9.0005
R867 iovss.n1824 iovss.n1739 9.0005
R868 iovss.n1790 iovss.n1739 9.0005
R869 iovss.n1827 iovss.n1739 9.0005
R870 iovss.n1789 iovss.n1739 9.0005
R871 iovss.n1830 iovss.n1739 9.0005
R872 iovss.n1788 iovss.n1739 9.0005
R873 iovss.n1832 iovss.n1739 9.0005
R874 iovss.n1787 iovss.n1739 9.0005
R875 iovss.n1835 iovss.n1739 9.0005
R876 iovss.n1786 iovss.n1739 9.0005
R877 iovss.n1837 iovss.n1739 9.0005
R878 iovss.n1785 iovss.n1739 9.0005
R879 iovss.n1840 iovss.n1739 9.0005
R880 iovss.n1784 iovss.n1739 9.0005
R881 iovss.n1841 iovss.n1739 9.0005
R882 iovss.n1870 iovss.n1739 9.0005
R883 iovss.n2290 iovss.n1739 9.0005
R884 iovss.n2292 iovss.n1723 9.0005
R885 iovss.n1801 iovss.n1723 9.0005
R886 iovss.n1799 iovss.n1723 9.0005
R887 iovss.n1804 iovss.n1723 9.0005
R888 iovss.n1798 iovss.n1723 9.0005
R889 iovss.n1807 iovss.n1723 9.0005
R890 iovss.n1797 iovss.n1723 9.0005
R891 iovss.n1809 iovss.n1723 9.0005
R892 iovss.n1796 iovss.n1723 9.0005
R893 iovss.n1812 iovss.n1723 9.0005
R894 iovss.n1795 iovss.n1723 9.0005
R895 iovss.n1814 iovss.n1723 9.0005
R896 iovss.n1794 iovss.n1723 9.0005
R897 iovss.n1817 iovss.n1723 9.0005
R898 iovss.n1793 iovss.n1723 9.0005
R899 iovss.n1819 iovss.n1723 9.0005
R900 iovss.n1792 iovss.n1723 9.0005
R901 iovss.n1822 iovss.n1723 9.0005
R902 iovss.n1791 iovss.n1723 9.0005
R903 iovss.n1824 iovss.n1723 9.0005
R904 iovss.n1790 iovss.n1723 9.0005
R905 iovss.n1827 iovss.n1723 9.0005
R906 iovss.n1789 iovss.n1723 9.0005
R907 iovss.n1830 iovss.n1723 9.0005
R908 iovss.n1788 iovss.n1723 9.0005
R909 iovss.n1832 iovss.n1723 9.0005
R910 iovss.n1787 iovss.n1723 9.0005
R911 iovss.n1835 iovss.n1723 9.0005
R912 iovss.n1786 iovss.n1723 9.0005
R913 iovss.n1837 iovss.n1723 9.0005
R914 iovss.n1785 iovss.n1723 9.0005
R915 iovss.n1840 iovss.n1723 9.0005
R916 iovss.n1784 iovss.n1723 9.0005
R917 iovss.n1841 iovss.n1723 9.0005
R918 iovss.n1870 iovss.n1723 9.0005
R919 iovss.n2290 iovss.n1723 9.0005
R920 iovss.n2292 iovss.n1740 9.0005
R921 iovss.n1801 iovss.n1740 9.0005
R922 iovss.n1799 iovss.n1740 9.0005
R923 iovss.n1804 iovss.n1740 9.0005
R924 iovss.n1798 iovss.n1740 9.0005
R925 iovss.n1807 iovss.n1740 9.0005
R926 iovss.n1797 iovss.n1740 9.0005
R927 iovss.n1809 iovss.n1740 9.0005
R928 iovss.n1796 iovss.n1740 9.0005
R929 iovss.n1812 iovss.n1740 9.0005
R930 iovss.n1795 iovss.n1740 9.0005
R931 iovss.n1814 iovss.n1740 9.0005
R932 iovss.n1794 iovss.n1740 9.0005
R933 iovss.n1817 iovss.n1740 9.0005
R934 iovss.n1793 iovss.n1740 9.0005
R935 iovss.n1819 iovss.n1740 9.0005
R936 iovss.n1792 iovss.n1740 9.0005
R937 iovss.n1822 iovss.n1740 9.0005
R938 iovss.n1791 iovss.n1740 9.0005
R939 iovss.n1824 iovss.n1740 9.0005
R940 iovss.n1790 iovss.n1740 9.0005
R941 iovss.n1827 iovss.n1740 9.0005
R942 iovss.n1789 iovss.n1740 9.0005
R943 iovss.n1830 iovss.n1740 9.0005
R944 iovss.n1788 iovss.n1740 9.0005
R945 iovss.n1832 iovss.n1740 9.0005
R946 iovss.n1787 iovss.n1740 9.0005
R947 iovss.n1835 iovss.n1740 9.0005
R948 iovss.n1786 iovss.n1740 9.0005
R949 iovss.n1837 iovss.n1740 9.0005
R950 iovss.n1785 iovss.n1740 9.0005
R951 iovss.n1840 iovss.n1740 9.0005
R952 iovss.n1784 iovss.n1740 9.0005
R953 iovss.n1841 iovss.n1740 9.0005
R954 iovss.n1870 iovss.n1740 9.0005
R955 iovss.n2290 iovss.n1740 9.0005
R956 iovss.n2292 iovss.n1722 9.0005
R957 iovss.n1801 iovss.n1722 9.0005
R958 iovss.n1799 iovss.n1722 9.0005
R959 iovss.n1804 iovss.n1722 9.0005
R960 iovss.n1798 iovss.n1722 9.0005
R961 iovss.n1807 iovss.n1722 9.0005
R962 iovss.n1797 iovss.n1722 9.0005
R963 iovss.n1809 iovss.n1722 9.0005
R964 iovss.n1796 iovss.n1722 9.0005
R965 iovss.n1812 iovss.n1722 9.0005
R966 iovss.n1795 iovss.n1722 9.0005
R967 iovss.n1814 iovss.n1722 9.0005
R968 iovss.n1794 iovss.n1722 9.0005
R969 iovss.n1817 iovss.n1722 9.0005
R970 iovss.n1793 iovss.n1722 9.0005
R971 iovss.n1819 iovss.n1722 9.0005
R972 iovss.n1792 iovss.n1722 9.0005
R973 iovss.n1822 iovss.n1722 9.0005
R974 iovss.n1791 iovss.n1722 9.0005
R975 iovss.n1824 iovss.n1722 9.0005
R976 iovss.n1790 iovss.n1722 9.0005
R977 iovss.n1827 iovss.n1722 9.0005
R978 iovss.n1789 iovss.n1722 9.0005
R979 iovss.n1830 iovss.n1722 9.0005
R980 iovss.n1788 iovss.n1722 9.0005
R981 iovss.n1832 iovss.n1722 9.0005
R982 iovss.n1787 iovss.n1722 9.0005
R983 iovss.n1835 iovss.n1722 9.0005
R984 iovss.n1786 iovss.n1722 9.0005
R985 iovss.n1837 iovss.n1722 9.0005
R986 iovss.n1785 iovss.n1722 9.0005
R987 iovss.n1840 iovss.n1722 9.0005
R988 iovss.n1784 iovss.n1722 9.0005
R989 iovss.n1841 iovss.n1722 9.0005
R990 iovss.n1870 iovss.n1722 9.0005
R991 iovss.n2290 iovss.n1722 9.0005
R992 iovss.n2292 iovss.n1741 9.0005
R993 iovss.n1801 iovss.n1741 9.0005
R994 iovss.n1799 iovss.n1741 9.0005
R995 iovss.n1804 iovss.n1741 9.0005
R996 iovss.n1798 iovss.n1741 9.0005
R997 iovss.n1807 iovss.n1741 9.0005
R998 iovss.n1797 iovss.n1741 9.0005
R999 iovss.n1809 iovss.n1741 9.0005
R1000 iovss.n1796 iovss.n1741 9.0005
R1001 iovss.n1812 iovss.n1741 9.0005
R1002 iovss.n1795 iovss.n1741 9.0005
R1003 iovss.n1814 iovss.n1741 9.0005
R1004 iovss.n1794 iovss.n1741 9.0005
R1005 iovss.n1817 iovss.n1741 9.0005
R1006 iovss.n1793 iovss.n1741 9.0005
R1007 iovss.n1819 iovss.n1741 9.0005
R1008 iovss.n1792 iovss.n1741 9.0005
R1009 iovss.n1822 iovss.n1741 9.0005
R1010 iovss.n1791 iovss.n1741 9.0005
R1011 iovss.n1824 iovss.n1741 9.0005
R1012 iovss.n1790 iovss.n1741 9.0005
R1013 iovss.n1827 iovss.n1741 9.0005
R1014 iovss.n1789 iovss.n1741 9.0005
R1015 iovss.n1830 iovss.n1741 9.0005
R1016 iovss.n1788 iovss.n1741 9.0005
R1017 iovss.n1832 iovss.n1741 9.0005
R1018 iovss.n1787 iovss.n1741 9.0005
R1019 iovss.n1835 iovss.n1741 9.0005
R1020 iovss.n1786 iovss.n1741 9.0005
R1021 iovss.n1837 iovss.n1741 9.0005
R1022 iovss.n1785 iovss.n1741 9.0005
R1023 iovss.n1840 iovss.n1741 9.0005
R1024 iovss.n1784 iovss.n1741 9.0005
R1025 iovss.n1841 iovss.n1741 9.0005
R1026 iovss.n1870 iovss.n1741 9.0005
R1027 iovss.n2290 iovss.n1741 9.0005
R1028 iovss.n2292 iovss.n1721 9.0005
R1029 iovss.n1801 iovss.n1721 9.0005
R1030 iovss.n1799 iovss.n1721 9.0005
R1031 iovss.n1804 iovss.n1721 9.0005
R1032 iovss.n1798 iovss.n1721 9.0005
R1033 iovss.n1807 iovss.n1721 9.0005
R1034 iovss.n1797 iovss.n1721 9.0005
R1035 iovss.n1809 iovss.n1721 9.0005
R1036 iovss.n1796 iovss.n1721 9.0005
R1037 iovss.n1812 iovss.n1721 9.0005
R1038 iovss.n1795 iovss.n1721 9.0005
R1039 iovss.n1814 iovss.n1721 9.0005
R1040 iovss.n1794 iovss.n1721 9.0005
R1041 iovss.n1817 iovss.n1721 9.0005
R1042 iovss.n1793 iovss.n1721 9.0005
R1043 iovss.n1819 iovss.n1721 9.0005
R1044 iovss.n1792 iovss.n1721 9.0005
R1045 iovss.n1822 iovss.n1721 9.0005
R1046 iovss.n1791 iovss.n1721 9.0005
R1047 iovss.n1824 iovss.n1721 9.0005
R1048 iovss.n1790 iovss.n1721 9.0005
R1049 iovss.n1827 iovss.n1721 9.0005
R1050 iovss.n1789 iovss.n1721 9.0005
R1051 iovss.n1830 iovss.n1721 9.0005
R1052 iovss.n1788 iovss.n1721 9.0005
R1053 iovss.n1832 iovss.n1721 9.0005
R1054 iovss.n1787 iovss.n1721 9.0005
R1055 iovss.n1835 iovss.n1721 9.0005
R1056 iovss.n1786 iovss.n1721 9.0005
R1057 iovss.n1837 iovss.n1721 9.0005
R1058 iovss.n1785 iovss.n1721 9.0005
R1059 iovss.n1840 iovss.n1721 9.0005
R1060 iovss.n1784 iovss.n1721 9.0005
R1061 iovss.n1841 iovss.n1721 9.0005
R1062 iovss.n1870 iovss.n1721 9.0005
R1063 iovss.n2290 iovss.n1721 9.0005
R1064 iovss.n2292 iovss.n1742 9.0005
R1065 iovss.n1801 iovss.n1742 9.0005
R1066 iovss.n1799 iovss.n1742 9.0005
R1067 iovss.n1804 iovss.n1742 9.0005
R1068 iovss.n1798 iovss.n1742 9.0005
R1069 iovss.n1807 iovss.n1742 9.0005
R1070 iovss.n1797 iovss.n1742 9.0005
R1071 iovss.n1809 iovss.n1742 9.0005
R1072 iovss.n1796 iovss.n1742 9.0005
R1073 iovss.n1812 iovss.n1742 9.0005
R1074 iovss.n1795 iovss.n1742 9.0005
R1075 iovss.n1814 iovss.n1742 9.0005
R1076 iovss.n1794 iovss.n1742 9.0005
R1077 iovss.n1817 iovss.n1742 9.0005
R1078 iovss.n1793 iovss.n1742 9.0005
R1079 iovss.n1819 iovss.n1742 9.0005
R1080 iovss.n1792 iovss.n1742 9.0005
R1081 iovss.n1822 iovss.n1742 9.0005
R1082 iovss.n1791 iovss.n1742 9.0005
R1083 iovss.n1824 iovss.n1742 9.0005
R1084 iovss.n1790 iovss.n1742 9.0005
R1085 iovss.n1827 iovss.n1742 9.0005
R1086 iovss.n1789 iovss.n1742 9.0005
R1087 iovss.n1830 iovss.n1742 9.0005
R1088 iovss.n1788 iovss.n1742 9.0005
R1089 iovss.n1832 iovss.n1742 9.0005
R1090 iovss.n1787 iovss.n1742 9.0005
R1091 iovss.n1835 iovss.n1742 9.0005
R1092 iovss.n1786 iovss.n1742 9.0005
R1093 iovss.n1837 iovss.n1742 9.0005
R1094 iovss.n1785 iovss.n1742 9.0005
R1095 iovss.n1840 iovss.n1742 9.0005
R1096 iovss.n1784 iovss.n1742 9.0005
R1097 iovss.n1841 iovss.n1742 9.0005
R1098 iovss.n1870 iovss.n1742 9.0005
R1099 iovss.n2290 iovss.n1742 9.0005
R1100 iovss.n2292 iovss.n1720 9.0005
R1101 iovss.n1801 iovss.n1720 9.0005
R1102 iovss.n1799 iovss.n1720 9.0005
R1103 iovss.n1804 iovss.n1720 9.0005
R1104 iovss.n1798 iovss.n1720 9.0005
R1105 iovss.n1807 iovss.n1720 9.0005
R1106 iovss.n1797 iovss.n1720 9.0005
R1107 iovss.n1809 iovss.n1720 9.0005
R1108 iovss.n1796 iovss.n1720 9.0005
R1109 iovss.n1812 iovss.n1720 9.0005
R1110 iovss.n1795 iovss.n1720 9.0005
R1111 iovss.n1814 iovss.n1720 9.0005
R1112 iovss.n1794 iovss.n1720 9.0005
R1113 iovss.n1817 iovss.n1720 9.0005
R1114 iovss.n1793 iovss.n1720 9.0005
R1115 iovss.n1819 iovss.n1720 9.0005
R1116 iovss.n1792 iovss.n1720 9.0005
R1117 iovss.n1822 iovss.n1720 9.0005
R1118 iovss.n1791 iovss.n1720 9.0005
R1119 iovss.n1824 iovss.n1720 9.0005
R1120 iovss.n1790 iovss.n1720 9.0005
R1121 iovss.n1827 iovss.n1720 9.0005
R1122 iovss.n1789 iovss.n1720 9.0005
R1123 iovss.n1830 iovss.n1720 9.0005
R1124 iovss.n1788 iovss.n1720 9.0005
R1125 iovss.n1832 iovss.n1720 9.0005
R1126 iovss.n1787 iovss.n1720 9.0005
R1127 iovss.n1835 iovss.n1720 9.0005
R1128 iovss.n1786 iovss.n1720 9.0005
R1129 iovss.n1837 iovss.n1720 9.0005
R1130 iovss.n1785 iovss.n1720 9.0005
R1131 iovss.n1840 iovss.n1720 9.0005
R1132 iovss.n1784 iovss.n1720 9.0005
R1133 iovss.n1841 iovss.n1720 9.0005
R1134 iovss.n1870 iovss.n1720 9.0005
R1135 iovss.n2290 iovss.n1720 9.0005
R1136 iovss.n2292 iovss.n1743 9.0005
R1137 iovss.n1801 iovss.n1743 9.0005
R1138 iovss.n1799 iovss.n1743 9.0005
R1139 iovss.n1804 iovss.n1743 9.0005
R1140 iovss.n1798 iovss.n1743 9.0005
R1141 iovss.n1807 iovss.n1743 9.0005
R1142 iovss.n1797 iovss.n1743 9.0005
R1143 iovss.n1809 iovss.n1743 9.0005
R1144 iovss.n1796 iovss.n1743 9.0005
R1145 iovss.n1812 iovss.n1743 9.0005
R1146 iovss.n1795 iovss.n1743 9.0005
R1147 iovss.n1814 iovss.n1743 9.0005
R1148 iovss.n1794 iovss.n1743 9.0005
R1149 iovss.n1817 iovss.n1743 9.0005
R1150 iovss.n1793 iovss.n1743 9.0005
R1151 iovss.n1819 iovss.n1743 9.0005
R1152 iovss.n1792 iovss.n1743 9.0005
R1153 iovss.n1822 iovss.n1743 9.0005
R1154 iovss.n1791 iovss.n1743 9.0005
R1155 iovss.n1824 iovss.n1743 9.0005
R1156 iovss.n1790 iovss.n1743 9.0005
R1157 iovss.n1827 iovss.n1743 9.0005
R1158 iovss.n1789 iovss.n1743 9.0005
R1159 iovss.n1830 iovss.n1743 9.0005
R1160 iovss.n1788 iovss.n1743 9.0005
R1161 iovss.n1832 iovss.n1743 9.0005
R1162 iovss.n1787 iovss.n1743 9.0005
R1163 iovss.n1835 iovss.n1743 9.0005
R1164 iovss.n1786 iovss.n1743 9.0005
R1165 iovss.n1837 iovss.n1743 9.0005
R1166 iovss.n1785 iovss.n1743 9.0005
R1167 iovss.n1840 iovss.n1743 9.0005
R1168 iovss.n1784 iovss.n1743 9.0005
R1169 iovss.n1841 iovss.n1743 9.0005
R1170 iovss.n1870 iovss.n1743 9.0005
R1171 iovss.n2290 iovss.n1743 9.0005
R1172 iovss.n2292 iovss.n1719 9.0005
R1173 iovss.n1801 iovss.n1719 9.0005
R1174 iovss.n1799 iovss.n1719 9.0005
R1175 iovss.n1804 iovss.n1719 9.0005
R1176 iovss.n1798 iovss.n1719 9.0005
R1177 iovss.n1807 iovss.n1719 9.0005
R1178 iovss.n1797 iovss.n1719 9.0005
R1179 iovss.n1809 iovss.n1719 9.0005
R1180 iovss.n1796 iovss.n1719 9.0005
R1181 iovss.n1812 iovss.n1719 9.0005
R1182 iovss.n1795 iovss.n1719 9.0005
R1183 iovss.n1814 iovss.n1719 9.0005
R1184 iovss.n1794 iovss.n1719 9.0005
R1185 iovss.n1817 iovss.n1719 9.0005
R1186 iovss.n1793 iovss.n1719 9.0005
R1187 iovss.n1819 iovss.n1719 9.0005
R1188 iovss.n1792 iovss.n1719 9.0005
R1189 iovss.n1822 iovss.n1719 9.0005
R1190 iovss.n1791 iovss.n1719 9.0005
R1191 iovss.n1824 iovss.n1719 9.0005
R1192 iovss.n1790 iovss.n1719 9.0005
R1193 iovss.n1827 iovss.n1719 9.0005
R1194 iovss.n1789 iovss.n1719 9.0005
R1195 iovss.n1830 iovss.n1719 9.0005
R1196 iovss.n1788 iovss.n1719 9.0005
R1197 iovss.n1832 iovss.n1719 9.0005
R1198 iovss.n1787 iovss.n1719 9.0005
R1199 iovss.n1835 iovss.n1719 9.0005
R1200 iovss.n1786 iovss.n1719 9.0005
R1201 iovss.n1837 iovss.n1719 9.0005
R1202 iovss.n1785 iovss.n1719 9.0005
R1203 iovss.n1840 iovss.n1719 9.0005
R1204 iovss.n1784 iovss.n1719 9.0005
R1205 iovss.n1841 iovss.n1719 9.0005
R1206 iovss.n1870 iovss.n1719 9.0005
R1207 iovss.n2290 iovss.n1719 9.0005
R1208 iovss.n2292 iovss.n1744 9.0005
R1209 iovss.n1801 iovss.n1744 9.0005
R1210 iovss.n1799 iovss.n1744 9.0005
R1211 iovss.n1804 iovss.n1744 9.0005
R1212 iovss.n1798 iovss.n1744 9.0005
R1213 iovss.n1807 iovss.n1744 9.0005
R1214 iovss.n1797 iovss.n1744 9.0005
R1215 iovss.n1809 iovss.n1744 9.0005
R1216 iovss.n1796 iovss.n1744 9.0005
R1217 iovss.n1812 iovss.n1744 9.0005
R1218 iovss.n1795 iovss.n1744 9.0005
R1219 iovss.n1814 iovss.n1744 9.0005
R1220 iovss.n1794 iovss.n1744 9.0005
R1221 iovss.n1817 iovss.n1744 9.0005
R1222 iovss.n1793 iovss.n1744 9.0005
R1223 iovss.n1819 iovss.n1744 9.0005
R1224 iovss.n1792 iovss.n1744 9.0005
R1225 iovss.n1822 iovss.n1744 9.0005
R1226 iovss.n1791 iovss.n1744 9.0005
R1227 iovss.n1824 iovss.n1744 9.0005
R1228 iovss.n1790 iovss.n1744 9.0005
R1229 iovss.n1827 iovss.n1744 9.0005
R1230 iovss.n1789 iovss.n1744 9.0005
R1231 iovss.n1830 iovss.n1744 9.0005
R1232 iovss.n1788 iovss.n1744 9.0005
R1233 iovss.n1832 iovss.n1744 9.0005
R1234 iovss.n1787 iovss.n1744 9.0005
R1235 iovss.n1835 iovss.n1744 9.0005
R1236 iovss.n1786 iovss.n1744 9.0005
R1237 iovss.n1837 iovss.n1744 9.0005
R1238 iovss.n1785 iovss.n1744 9.0005
R1239 iovss.n1840 iovss.n1744 9.0005
R1240 iovss.n1784 iovss.n1744 9.0005
R1241 iovss.n1841 iovss.n1744 9.0005
R1242 iovss.n1870 iovss.n1744 9.0005
R1243 iovss.n2290 iovss.n1744 9.0005
R1244 iovss.n2292 iovss.n1718 9.0005
R1245 iovss.n1801 iovss.n1718 9.0005
R1246 iovss.n1799 iovss.n1718 9.0005
R1247 iovss.n1804 iovss.n1718 9.0005
R1248 iovss.n1798 iovss.n1718 9.0005
R1249 iovss.n1807 iovss.n1718 9.0005
R1250 iovss.n1797 iovss.n1718 9.0005
R1251 iovss.n1809 iovss.n1718 9.0005
R1252 iovss.n1796 iovss.n1718 9.0005
R1253 iovss.n1812 iovss.n1718 9.0005
R1254 iovss.n1795 iovss.n1718 9.0005
R1255 iovss.n1814 iovss.n1718 9.0005
R1256 iovss.n1794 iovss.n1718 9.0005
R1257 iovss.n1817 iovss.n1718 9.0005
R1258 iovss.n1793 iovss.n1718 9.0005
R1259 iovss.n1819 iovss.n1718 9.0005
R1260 iovss.n1792 iovss.n1718 9.0005
R1261 iovss.n1822 iovss.n1718 9.0005
R1262 iovss.n1791 iovss.n1718 9.0005
R1263 iovss.n1824 iovss.n1718 9.0005
R1264 iovss.n1790 iovss.n1718 9.0005
R1265 iovss.n1827 iovss.n1718 9.0005
R1266 iovss.n1789 iovss.n1718 9.0005
R1267 iovss.n1830 iovss.n1718 9.0005
R1268 iovss.n1788 iovss.n1718 9.0005
R1269 iovss.n1832 iovss.n1718 9.0005
R1270 iovss.n1787 iovss.n1718 9.0005
R1271 iovss.n1835 iovss.n1718 9.0005
R1272 iovss.n1786 iovss.n1718 9.0005
R1273 iovss.n1837 iovss.n1718 9.0005
R1274 iovss.n1785 iovss.n1718 9.0005
R1275 iovss.n1840 iovss.n1718 9.0005
R1276 iovss.n1784 iovss.n1718 9.0005
R1277 iovss.n1841 iovss.n1718 9.0005
R1278 iovss.n1870 iovss.n1718 9.0005
R1279 iovss.n2290 iovss.n1718 9.0005
R1280 iovss.n2292 iovss.n1745 9.0005
R1281 iovss.n1801 iovss.n1745 9.0005
R1282 iovss.n1799 iovss.n1745 9.0005
R1283 iovss.n1804 iovss.n1745 9.0005
R1284 iovss.n1798 iovss.n1745 9.0005
R1285 iovss.n1807 iovss.n1745 9.0005
R1286 iovss.n1797 iovss.n1745 9.0005
R1287 iovss.n1809 iovss.n1745 9.0005
R1288 iovss.n1796 iovss.n1745 9.0005
R1289 iovss.n1812 iovss.n1745 9.0005
R1290 iovss.n1795 iovss.n1745 9.0005
R1291 iovss.n1814 iovss.n1745 9.0005
R1292 iovss.n1794 iovss.n1745 9.0005
R1293 iovss.n1817 iovss.n1745 9.0005
R1294 iovss.n1793 iovss.n1745 9.0005
R1295 iovss.n1819 iovss.n1745 9.0005
R1296 iovss.n1792 iovss.n1745 9.0005
R1297 iovss.n1822 iovss.n1745 9.0005
R1298 iovss.n1791 iovss.n1745 9.0005
R1299 iovss.n1824 iovss.n1745 9.0005
R1300 iovss.n1790 iovss.n1745 9.0005
R1301 iovss.n1827 iovss.n1745 9.0005
R1302 iovss.n1789 iovss.n1745 9.0005
R1303 iovss.n1830 iovss.n1745 9.0005
R1304 iovss.n1788 iovss.n1745 9.0005
R1305 iovss.n1832 iovss.n1745 9.0005
R1306 iovss.n1787 iovss.n1745 9.0005
R1307 iovss.n1835 iovss.n1745 9.0005
R1308 iovss.n1786 iovss.n1745 9.0005
R1309 iovss.n1837 iovss.n1745 9.0005
R1310 iovss.n1785 iovss.n1745 9.0005
R1311 iovss.n1840 iovss.n1745 9.0005
R1312 iovss.n1784 iovss.n1745 9.0005
R1313 iovss.n1841 iovss.n1745 9.0005
R1314 iovss.n1870 iovss.n1745 9.0005
R1315 iovss.n2290 iovss.n1745 9.0005
R1316 iovss.n2292 iovss.n1717 9.0005
R1317 iovss.n1801 iovss.n1717 9.0005
R1318 iovss.n1799 iovss.n1717 9.0005
R1319 iovss.n1804 iovss.n1717 9.0005
R1320 iovss.n1798 iovss.n1717 9.0005
R1321 iovss.n1807 iovss.n1717 9.0005
R1322 iovss.n1797 iovss.n1717 9.0005
R1323 iovss.n1809 iovss.n1717 9.0005
R1324 iovss.n1796 iovss.n1717 9.0005
R1325 iovss.n1812 iovss.n1717 9.0005
R1326 iovss.n1795 iovss.n1717 9.0005
R1327 iovss.n1814 iovss.n1717 9.0005
R1328 iovss.n1794 iovss.n1717 9.0005
R1329 iovss.n1817 iovss.n1717 9.0005
R1330 iovss.n1793 iovss.n1717 9.0005
R1331 iovss.n1819 iovss.n1717 9.0005
R1332 iovss.n1792 iovss.n1717 9.0005
R1333 iovss.n1822 iovss.n1717 9.0005
R1334 iovss.n1791 iovss.n1717 9.0005
R1335 iovss.n1824 iovss.n1717 9.0005
R1336 iovss.n1790 iovss.n1717 9.0005
R1337 iovss.n1827 iovss.n1717 9.0005
R1338 iovss.n1789 iovss.n1717 9.0005
R1339 iovss.n1830 iovss.n1717 9.0005
R1340 iovss.n1788 iovss.n1717 9.0005
R1341 iovss.n1832 iovss.n1717 9.0005
R1342 iovss.n1787 iovss.n1717 9.0005
R1343 iovss.n1835 iovss.n1717 9.0005
R1344 iovss.n1786 iovss.n1717 9.0005
R1345 iovss.n1837 iovss.n1717 9.0005
R1346 iovss.n1785 iovss.n1717 9.0005
R1347 iovss.n1840 iovss.n1717 9.0005
R1348 iovss.n1784 iovss.n1717 9.0005
R1349 iovss.n1841 iovss.n1717 9.0005
R1350 iovss.n1870 iovss.n1717 9.0005
R1351 iovss.n2290 iovss.n1717 9.0005
R1352 iovss.n2292 iovss.n1746 9.0005
R1353 iovss.n1801 iovss.n1746 9.0005
R1354 iovss.n1799 iovss.n1746 9.0005
R1355 iovss.n1804 iovss.n1746 9.0005
R1356 iovss.n1798 iovss.n1746 9.0005
R1357 iovss.n1807 iovss.n1746 9.0005
R1358 iovss.n1797 iovss.n1746 9.0005
R1359 iovss.n1809 iovss.n1746 9.0005
R1360 iovss.n1796 iovss.n1746 9.0005
R1361 iovss.n1812 iovss.n1746 9.0005
R1362 iovss.n1795 iovss.n1746 9.0005
R1363 iovss.n1814 iovss.n1746 9.0005
R1364 iovss.n1794 iovss.n1746 9.0005
R1365 iovss.n1817 iovss.n1746 9.0005
R1366 iovss.n1793 iovss.n1746 9.0005
R1367 iovss.n1819 iovss.n1746 9.0005
R1368 iovss.n1792 iovss.n1746 9.0005
R1369 iovss.n1822 iovss.n1746 9.0005
R1370 iovss.n1791 iovss.n1746 9.0005
R1371 iovss.n1824 iovss.n1746 9.0005
R1372 iovss.n1790 iovss.n1746 9.0005
R1373 iovss.n1827 iovss.n1746 9.0005
R1374 iovss.n1789 iovss.n1746 9.0005
R1375 iovss.n1830 iovss.n1746 9.0005
R1376 iovss.n1788 iovss.n1746 9.0005
R1377 iovss.n1832 iovss.n1746 9.0005
R1378 iovss.n1787 iovss.n1746 9.0005
R1379 iovss.n1835 iovss.n1746 9.0005
R1380 iovss.n1786 iovss.n1746 9.0005
R1381 iovss.n1837 iovss.n1746 9.0005
R1382 iovss.n1785 iovss.n1746 9.0005
R1383 iovss.n1840 iovss.n1746 9.0005
R1384 iovss.n1784 iovss.n1746 9.0005
R1385 iovss.n1841 iovss.n1746 9.0005
R1386 iovss.n1870 iovss.n1746 9.0005
R1387 iovss.n2290 iovss.n1746 9.0005
R1388 iovss.n2292 iovss.n1716 9.0005
R1389 iovss.n1801 iovss.n1716 9.0005
R1390 iovss.n1799 iovss.n1716 9.0005
R1391 iovss.n1804 iovss.n1716 9.0005
R1392 iovss.n1798 iovss.n1716 9.0005
R1393 iovss.n1807 iovss.n1716 9.0005
R1394 iovss.n1797 iovss.n1716 9.0005
R1395 iovss.n1809 iovss.n1716 9.0005
R1396 iovss.n1796 iovss.n1716 9.0005
R1397 iovss.n1812 iovss.n1716 9.0005
R1398 iovss.n1795 iovss.n1716 9.0005
R1399 iovss.n1814 iovss.n1716 9.0005
R1400 iovss.n1794 iovss.n1716 9.0005
R1401 iovss.n1817 iovss.n1716 9.0005
R1402 iovss.n1793 iovss.n1716 9.0005
R1403 iovss.n1819 iovss.n1716 9.0005
R1404 iovss.n1792 iovss.n1716 9.0005
R1405 iovss.n1822 iovss.n1716 9.0005
R1406 iovss.n1791 iovss.n1716 9.0005
R1407 iovss.n1824 iovss.n1716 9.0005
R1408 iovss.n1790 iovss.n1716 9.0005
R1409 iovss.n1827 iovss.n1716 9.0005
R1410 iovss.n1789 iovss.n1716 9.0005
R1411 iovss.n1830 iovss.n1716 9.0005
R1412 iovss.n1788 iovss.n1716 9.0005
R1413 iovss.n1832 iovss.n1716 9.0005
R1414 iovss.n1787 iovss.n1716 9.0005
R1415 iovss.n1835 iovss.n1716 9.0005
R1416 iovss.n1786 iovss.n1716 9.0005
R1417 iovss.n1837 iovss.n1716 9.0005
R1418 iovss.n1785 iovss.n1716 9.0005
R1419 iovss.n1840 iovss.n1716 9.0005
R1420 iovss.n1784 iovss.n1716 9.0005
R1421 iovss.n1841 iovss.n1716 9.0005
R1422 iovss.n1870 iovss.n1716 9.0005
R1423 iovss.n2290 iovss.n1716 9.0005
R1424 iovss.n2292 iovss.n1747 9.0005
R1425 iovss.n1801 iovss.n1747 9.0005
R1426 iovss.n1799 iovss.n1747 9.0005
R1427 iovss.n1804 iovss.n1747 9.0005
R1428 iovss.n1798 iovss.n1747 9.0005
R1429 iovss.n1807 iovss.n1747 9.0005
R1430 iovss.n1797 iovss.n1747 9.0005
R1431 iovss.n1809 iovss.n1747 9.0005
R1432 iovss.n1796 iovss.n1747 9.0005
R1433 iovss.n1812 iovss.n1747 9.0005
R1434 iovss.n1795 iovss.n1747 9.0005
R1435 iovss.n1814 iovss.n1747 9.0005
R1436 iovss.n1794 iovss.n1747 9.0005
R1437 iovss.n1817 iovss.n1747 9.0005
R1438 iovss.n1793 iovss.n1747 9.0005
R1439 iovss.n1819 iovss.n1747 9.0005
R1440 iovss.n1792 iovss.n1747 9.0005
R1441 iovss.n1822 iovss.n1747 9.0005
R1442 iovss.n1791 iovss.n1747 9.0005
R1443 iovss.n1824 iovss.n1747 9.0005
R1444 iovss.n1790 iovss.n1747 9.0005
R1445 iovss.n1827 iovss.n1747 9.0005
R1446 iovss.n1789 iovss.n1747 9.0005
R1447 iovss.n1830 iovss.n1747 9.0005
R1448 iovss.n1788 iovss.n1747 9.0005
R1449 iovss.n1832 iovss.n1747 9.0005
R1450 iovss.n1787 iovss.n1747 9.0005
R1451 iovss.n1835 iovss.n1747 9.0005
R1452 iovss.n1786 iovss.n1747 9.0005
R1453 iovss.n1837 iovss.n1747 9.0005
R1454 iovss.n1785 iovss.n1747 9.0005
R1455 iovss.n1840 iovss.n1747 9.0005
R1456 iovss.n1784 iovss.n1747 9.0005
R1457 iovss.n1841 iovss.n1747 9.0005
R1458 iovss.n1870 iovss.n1747 9.0005
R1459 iovss.n2290 iovss.n1747 9.0005
R1460 iovss.n2292 iovss.n1715 9.0005
R1461 iovss.n1801 iovss.n1715 9.0005
R1462 iovss.n1799 iovss.n1715 9.0005
R1463 iovss.n1804 iovss.n1715 9.0005
R1464 iovss.n1798 iovss.n1715 9.0005
R1465 iovss.n1807 iovss.n1715 9.0005
R1466 iovss.n1797 iovss.n1715 9.0005
R1467 iovss.n1809 iovss.n1715 9.0005
R1468 iovss.n1796 iovss.n1715 9.0005
R1469 iovss.n1812 iovss.n1715 9.0005
R1470 iovss.n1795 iovss.n1715 9.0005
R1471 iovss.n1814 iovss.n1715 9.0005
R1472 iovss.n1794 iovss.n1715 9.0005
R1473 iovss.n1817 iovss.n1715 9.0005
R1474 iovss.n1793 iovss.n1715 9.0005
R1475 iovss.n1819 iovss.n1715 9.0005
R1476 iovss.n1792 iovss.n1715 9.0005
R1477 iovss.n1822 iovss.n1715 9.0005
R1478 iovss.n1791 iovss.n1715 9.0005
R1479 iovss.n1824 iovss.n1715 9.0005
R1480 iovss.n1790 iovss.n1715 9.0005
R1481 iovss.n1827 iovss.n1715 9.0005
R1482 iovss.n1789 iovss.n1715 9.0005
R1483 iovss.n1830 iovss.n1715 9.0005
R1484 iovss.n1788 iovss.n1715 9.0005
R1485 iovss.n1832 iovss.n1715 9.0005
R1486 iovss.n1787 iovss.n1715 9.0005
R1487 iovss.n1835 iovss.n1715 9.0005
R1488 iovss.n1786 iovss.n1715 9.0005
R1489 iovss.n1837 iovss.n1715 9.0005
R1490 iovss.n1785 iovss.n1715 9.0005
R1491 iovss.n1840 iovss.n1715 9.0005
R1492 iovss.n1784 iovss.n1715 9.0005
R1493 iovss.n1841 iovss.n1715 9.0005
R1494 iovss.n1870 iovss.n1715 9.0005
R1495 iovss.n2290 iovss.n1715 9.0005
R1496 iovss.n2292 iovss.n1748 9.0005
R1497 iovss.n1801 iovss.n1748 9.0005
R1498 iovss.n1799 iovss.n1748 9.0005
R1499 iovss.n1804 iovss.n1748 9.0005
R1500 iovss.n1798 iovss.n1748 9.0005
R1501 iovss.n1807 iovss.n1748 9.0005
R1502 iovss.n1797 iovss.n1748 9.0005
R1503 iovss.n1809 iovss.n1748 9.0005
R1504 iovss.n1796 iovss.n1748 9.0005
R1505 iovss.n1812 iovss.n1748 9.0005
R1506 iovss.n1795 iovss.n1748 9.0005
R1507 iovss.n1814 iovss.n1748 9.0005
R1508 iovss.n1794 iovss.n1748 9.0005
R1509 iovss.n1817 iovss.n1748 9.0005
R1510 iovss.n1793 iovss.n1748 9.0005
R1511 iovss.n1819 iovss.n1748 9.0005
R1512 iovss.n1792 iovss.n1748 9.0005
R1513 iovss.n1822 iovss.n1748 9.0005
R1514 iovss.n1791 iovss.n1748 9.0005
R1515 iovss.n1824 iovss.n1748 9.0005
R1516 iovss.n1790 iovss.n1748 9.0005
R1517 iovss.n1827 iovss.n1748 9.0005
R1518 iovss.n1789 iovss.n1748 9.0005
R1519 iovss.n1830 iovss.n1748 9.0005
R1520 iovss.n1788 iovss.n1748 9.0005
R1521 iovss.n1832 iovss.n1748 9.0005
R1522 iovss.n1787 iovss.n1748 9.0005
R1523 iovss.n1835 iovss.n1748 9.0005
R1524 iovss.n1786 iovss.n1748 9.0005
R1525 iovss.n1837 iovss.n1748 9.0005
R1526 iovss.n1785 iovss.n1748 9.0005
R1527 iovss.n1840 iovss.n1748 9.0005
R1528 iovss.n1784 iovss.n1748 9.0005
R1529 iovss.n1841 iovss.n1748 9.0005
R1530 iovss.n1870 iovss.n1748 9.0005
R1531 iovss.n2290 iovss.n1748 9.0005
R1532 iovss.n2292 iovss.n1714 9.0005
R1533 iovss.n1801 iovss.n1714 9.0005
R1534 iovss.n1799 iovss.n1714 9.0005
R1535 iovss.n1804 iovss.n1714 9.0005
R1536 iovss.n1798 iovss.n1714 9.0005
R1537 iovss.n1807 iovss.n1714 9.0005
R1538 iovss.n1797 iovss.n1714 9.0005
R1539 iovss.n1809 iovss.n1714 9.0005
R1540 iovss.n1796 iovss.n1714 9.0005
R1541 iovss.n1812 iovss.n1714 9.0005
R1542 iovss.n1795 iovss.n1714 9.0005
R1543 iovss.n1814 iovss.n1714 9.0005
R1544 iovss.n1794 iovss.n1714 9.0005
R1545 iovss.n1817 iovss.n1714 9.0005
R1546 iovss.n1793 iovss.n1714 9.0005
R1547 iovss.n1819 iovss.n1714 9.0005
R1548 iovss.n1792 iovss.n1714 9.0005
R1549 iovss.n1822 iovss.n1714 9.0005
R1550 iovss.n1791 iovss.n1714 9.0005
R1551 iovss.n1824 iovss.n1714 9.0005
R1552 iovss.n1790 iovss.n1714 9.0005
R1553 iovss.n1827 iovss.n1714 9.0005
R1554 iovss.n1789 iovss.n1714 9.0005
R1555 iovss.n1830 iovss.n1714 9.0005
R1556 iovss.n1788 iovss.n1714 9.0005
R1557 iovss.n1832 iovss.n1714 9.0005
R1558 iovss.n1787 iovss.n1714 9.0005
R1559 iovss.n1835 iovss.n1714 9.0005
R1560 iovss.n1786 iovss.n1714 9.0005
R1561 iovss.n1837 iovss.n1714 9.0005
R1562 iovss.n1785 iovss.n1714 9.0005
R1563 iovss.n1840 iovss.n1714 9.0005
R1564 iovss.n1784 iovss.n1714 9.0005
R1565 iovss.n1841 iovss.n1714 9.0005
R1566 iovss.n1870 iovss.n1714 9.0005
R1567 iovss.n2290 iovss.n1714 9.0005
R1568 iovss.n2292 iovss.n1749 9.0005
R1569 iovss.n1801 iovss.n1749 9.0005
R1570 iovss.n1799 iovss.n1749 9.0005
R1571 iovss.n1804 iovss.n1749 9.0005
R1572 iovss.n1798 iovss.n1749 9.0005
R1573 iovss.n1807 iovss.n1749 9.0005
R1574 iovss.n1797 iovss.n1749 9.0005
R1575 iovss.n1809 iovss.n1749 9.0005
R1576 iovss.n1796 iovss.n1749 9.0005
R1577 iovss.n1812 iovss.n1749 9.0005
R1578 iovss.n1795 iovss.n1749 9.0005
R1579 iovss.n1814 iovss.n1749 9.0005
R1580 iovss.n1794 iovss.n1749 9.0005
R1581 iovss.n1817 iovss.n1749 9.0005
R1582 iovss.n1793 iovss.n1749 9.0005
R1583 iovss.n1819 iovss.n1749 9.0005
R1584 iovss.n1792 iovss.n1749 9.0005
R1585 iovss.n1822 iovss.n1749 9.0005
R1586 iovss.n1791 iovss.n1749 9.0005
R1587 iovss.n1824 iovss.n1749 9.0005
R1588 iovss.n1790 iovss.n1749 9.0005
R1589 iovss.n1827 iovss.n1749 9.0005
R1590 iovss.n1789 iovss.n1749 9.0005
R1591 iovss.n1830 iovss.n1749 9.0005
R1592 iovss.n1788 iovss.n1749 9.0005
R1593 iovss.n1832 iovss.n1749 9.0005
R1594 iovss.n1787 iovss.n1749 9.0005
R1595 iovss.n1835 iovss.n1749 9.0005
R1596 iovss.n1786 iovss.n1749 9.0005
R1597 iovss.n1837 iovss.n1749 9.0005
R1598 iovss.n1785 iovss.n1749 9.0005
R1599 iovss.n1840 iovss.n1749 9.0005
R1600 iovss.n1784 iovss.n1749 9.0005
R1601 iovss.n1841 iovss.n1749 9.0005
R1602 iovss.n1870 iovss.n1749 9.0005
R1603 iovss.n2290 iovss.n1749 9.0005
R1604 iovss.n2292 iovss.n1713 9.0005
R1605 iovss.n1801 iovss.n1713 9.0005
R1606 iovss.n1799 iovss.n1713 9.0005
R1607 iovss.n1804 iovss.n1713 9.0005
R1608 iovss.n1798 iovss.n1713 9.0005
R1609 iovss.n1807 iovss.n1713 9.0005
R1610 iovss.n1797 iovss.n1713 9.0005
R1611 iovss.n1809 iovss.n1713 9.0005
R1612 iovss.n1796 iovss.n1713 9.0005
R1613 iovss.n1812 iovss.n1713 9.0005
R1614 iovss.n1795 iovss.n1713 9.0005
R1615 iovss.n1814 iovss.n1713 9.0005
R1616 iovss.n1794 iovss.n1713 9.0005
R1617 iovss.n1817 iovss.n1713 9.0005
R1618 iovss.n1793 iovss.n1713 9.0005
R1619 iovss.n1819 iovss.n1713 9.0005
R1620 iovss.n1792 iovss.n1713 9.0005
R1621 iovss.n1822 iovss.n1713 9.0005
R1622 iovss.n1791 iovss.n1713 9.0005
R1623 iovss.n1824 iovss.n1713 9.0005
R1624 iovss.n1790 iovss.n1713 9.0005
R1625 iovss.n1827 iovss.n1713 9.0005
R1626 iovss.n1789 iovss.n1713 9.0005
R1627 iovss.n1830 iovss.n1713 9.0005
R1628 iovss.n1788 iovss.n1713 9.0005
R1629 iovss.n1832 iovss.n1713 9.0005
R1630 iovss.n1787 iovss.n1713 9.0005
R1631 iovss.n1835 iovss.n1713 9.0005
R1632 iovss.n1786 iovss.n1713 9.0005
R1633 iovss.n1837 iovss.n1713 9.0005
R1634 iovss.n1785 iovss.n1713 9.0005
R1635 iovss.n1840 iovss.n1713 9.0005
R1636 iovss.n1784 iovss.n1713 9.0005
R1637 iovss.n1841 iovss.n1713 9.0005
R1638 iovss.n1870 iovss.n1713 9.0005
R1639 iovss.n2290 iovss.n1713 9.0005
R1640 iovss.n2292 iovss.n1750 9.0005
R1641 iovss.n1801 iovss.n1750 9.0005
R1642 iovss.n1799 iovss.n1750 9.0005
R1643 iovss.n1804 iovss.n1750 9.0005
R1644 iovss.n1798 iovss.n1750 9.0005
R1645 iovss.n1807 iovss.n1750 9.0005
R1646 iovss.n1797 iovss.n1750 9.0005
R1647 iovss.n1809 iovss.n1750 9.0005
R1648 iovss.n1796 iovss.n1750 9.0005
R1649 iovss.n1812 iovss.n1750 9.0005
R1650 iovss.n1795 iovss.n1750 9.0005
R1651 iovss.n1814 iovss.n1750 9.0005
R1652 iovss.n1794 iovss.n1750 9.0005
R1653 iovss.n1817 iovss.n1750 9.0005
R1654 iovss.n1793 iovss.n1750 9.0005
R1655 iovss.n1819 iovss.n1750 9.0005
R1656 iovss.n1792 iovss.n1750 9.0005
R1657 iovss.n1822 iovss.n1750 9.0005
R1658 iovss.n1791 iovss.n1750 9.0005
R1659 iovss.n1824 iovss.n1750 9.0005
R1660 iovss.n1790 iovss.n1750 9.0005
R1661 iovss.n1827 iovss.n1750 9.0005
R1662 iovss.n1789 iovss.n1750 9.0005
R1663 iovss.n1830 iovss.n1750 9.0005
R1664 iovss.n1788 iovss.n1750 9.0005
R1665 iovss.n1832 iovss.n1750 9.0005
R1666 iovss.n1787 iovss.n1750 9.0005
R1667 iovss.n1835 iovss.n1750 9.0005
R1668 iovss.n1786 iovss.n1750 9.0005
R1669 iovss.n1837 iovss.n1750 9.0005
R1670 iovss.n1785 iovss.n1750 9.0005
R1671 iovss.n1840 iovss.n1750 9.0005
R1672 iovss.n1784 iovss.n1750 9.0005
R1673 iovss.n1841 iovss.n1750 9.0005
R1674 iovss.n1870 iovss.n1750 9.0005
R1675 iovss.n2290 iovss.n1750 9.0005
R1676 iovss.n2292 iovss.n1712 9.0005
R1677 iovss.n1801 iovss.n1712 9.0005
R1678 iovss.n1799 iovss.n1712 9.0005
R1679 iovss.n1804 iovss.n1712 9.0005
R1680 iovss.n1798 iovss.n1712 9.0005
R1681 iovss.n1807 iovss.n1712 9.0005
R1682 iovss.n1797 iovss.n1712 9.0005
R1683 iovss.n1809 iovss.n1712 9.0005
R1684 iovss.n1796 iovss.n1712 9.0005
R1685 iovss.n1812 iovss.n1712 9.0005
R1686 iovss.n1795 iovss.n1712 9.0005
R1687 iovss.n1814 iovss.n1712 9.0005
R1688 iovss.n1794 iovss.n1712 9.0005
R1689 iovss.n1817 iovss.n1712 9.0005
R1690 iovss.n1793 iovss.n1712 9.0005
R1691 iovss.n1819 iovss.n1712 9.0005
R1692 iovss.n1792 iovss.n1712 9.0005
R1693 iovss.n1822 iovss.n1712 9.0005
R1694 iovss.n1791 iovss.n1712 9.0005
R1695 iovss.n1824 iovss.n1712 9.0005
R1696 iovss.n1790 iovss.n1712 9.0005
R1697 iovss.n1827 iovss.n1712 9.0005
R1698 iovss.n1789 iovss.n1712 9.0005
R1699 iovss.n1830 iovss.n1712 9.0005
R1700 iovss.n1788 iovss.n1712 9.0005
R1701 iovss.n1832 iovss.n1712 9.0005
R1702 iovss.n1787 iovss.n1712 9.0005
R1703 iovss.n1835 iovss.n1712 9.0005
R1704 iovss.n1786 iovss.n1712 9.0005
R1705 iovss.n1837 iovss.n1712 9.0005
R1706 iovss.n1785 iovss.n1712 9.0005
R1707 iovss.n1840 iovss.n1712 9.0005
R1708 iovss.n1784 iovss.n1712 9.0005
R1709 iovss.n1841 iovss.n1712 9.0005
R1710 iovss.n1870 iovss.n1712 9.0005
R1711 iovss.n2290 iovss.n1712 9.0005
R1712 iovss.n2292 iovss.n1751 9.0005
R1713 iovss.n1801 iovss.n1751 9.0005
R1714 iovss.n1799 iovss.n1751 9.0005
R1715 iovss.n1804 iovss.n1751 9.0005
R1716 iovss.n1798 iovss.n1751 9.0005
R1717 iovss.n1807 iovss.n1751 9.0005
R1718 iovss.n1797 iovss.n1751 9.0005
R1719 iovss.n1809 iovss.n1751 9.0005
R1720 iovss.n1796 iovss.n1751 9.0005
R1721 iovss.n1812 iovss.n1751 9.0005
R1722 iovss.n1795 iovss.n1751 9.0005
R1723 iovss.n1814 iovss.n1751 9.0005
R1724 iovss.n1794 iovss.n1751 9.0005
R1725 iovss.n1817 iovss.n1751 9.0005
R1726 iovss.n1793 iovss.n1751 9.0005
R1727 iovss.n1819 iovss.n1751 9.0005
R1728 iovss.n1792 iovss.n1751 9.0005
R1729 iovss.n1822 iovss.n1751 9.0005
R1730 iovss.n1791 iovss.n1751 9.0005
R1731 iovss.n1824 iovss.n1751 9.0005
R1732 iovss.n1790 iovss.n1751 9.0005
R1733 iovss.n1827 iovss.n1751 9.0005
R1734 iovss.n1789 iovss.n1751 9.0005
R1735 iovss.n1830 iovss.n1751 9.0005
R1736 iovss.n1788 iovss.n1751 9.0005
R1737 iovss.n1832 iovss.n1751 9.0005
R1738 iovss.n1787 iovss.n1751 9.0005
R1739 iovss.n1835 iovss.n1751 9.0005
R1740 iovss.n1786 iovss.n1751 9.0005
R1741 iovss.n1837 iovss.n1751 9.0005
R1742 iovss.n1785 iovss.n1751 9.0005
R1743 iovss.n1840 iovss.n1751 9.0005
R1744 iovss.n1784 iovss.n1751 9.0005
R1745 iovss.n1841 iovss.n1751 9.0005
R1746 iovss.n1870 iovss.n1751 9.0005
R1747 iovss.n2290 iovss.n1751 9.0005
R1748 iovss.n2292 iovss.n1711 9.0005
R1749 iovss.n1801 iovss.n1711 9.0005
R1750 iovss.n1799 iovss.n1711 9.0005
R1751 iovss.n1804 iovss.n1711 9.0005
R1752 iovss.n1798 iovss.n1711 9.0005
R1753 iovss.n1807 iovss.n1711 9.0005
R1754 iovss.n1797 iovss.n1711 9.0005
R1755 iovss.n1809 iovss.n1711 9.0005
R1756 iovss.n1796 iovss.n1711 9.0005
R1757 iovss.n1812 iovss.n1711 9.0005
R1758 iovss.n1795 iovss.n1711 9.0005
R1759 iovss.n1814 iovss.n1711 9.0005
R1760 iovss.n1794 iovss.n1711 9.0005
R1761 iovss.n1817 iovss.n1711 9.0005
R1762 iovss.n1793 iovss.n1711 9.0005
R1763 iovss.n1819 iovss.n1711 9.0005
R1764 iovss.n1792 iovss.n1711 9.0005
R1765 iovss.n1822 iovss.n1711 9.0005
R1766 iovss.n1791 iovss.n1711 9.0005
R1767 iovss.n1824 iovss.n1711 9.0005
R1768 iovss.n1790 iovss.n1711 9.0005
R1769 iovss.n1827 iovss.n1711 9.0005
R1770 iovss.n1789 iovss.n1711 9.0005
R1771 iovss.n1830 iovss.n1711 9.0005
R1772 iovss.n1788 iovss.n1711 9.0005
R1773 iovss.n1832 iovss.n1711 9.0005
R1774 iovss.n1787 iovss.n1711 9.0005
R1775 iovss.n1835 iovss.n1711 9.0005
R1776 iovss.n1786 iovss.n1711 9.0005
R1777 iovss.n1837 iovss.n1711 9.0005
R1778 iovss.n1785 iovss.n1711 9.0005
R1779 iovss.n1840 iovss.n1711 9.0005
R1780 iovss.n1784 iovss.n1711 9.0005
R1781 iovss.n1841 iovss.n1711 9.0005
R1782 iovss.n1870 iovss.n1711 9.0005
R1783 iovss.n2290 iovss.n1711 9.0005
R1784 iovss.n2292 iovss.n1752 9.0005
R1785 iovss.n1801 iovss.n1752 9.0005
R1786 iovss.n1799 iovss.n1752 9.0005
R1787 iovss.n1804 iovss.n1752 9.0005
R1788 iovss.n1798 iovss.n1752 9.0005
R1789 iovss.n1807 iovss.n1752 9.0005
R1790 iovss.n1797 iovss.n1752 9.0005
R1791 iovss.n1809 iovss.n1752 9.0005
R1792 iovss.n1796 iovss.n1752 9.0005
R1793 iovss.n1812 iovss.n1752 9.0005
R1794 iovss.n1795 iovss.n1752 9.0005
R1795 iovss.n1814 iovss.n1752 9.0005
R1796 iovss.n1794 iovss.n1752 9.0005
R1797 iovss.n1817 iovss.n1752 9.0005
R1798 iovss.n1793 iovss.n1752 9.0005
R1799 iovss.n1819 iovss.n1752 9.0005
R1800 iovss.n1792 iovss.n1752 9.0005
R1801 iovss.n1822 iovss.n1752 9.0005
R1802 iovss.n1791 iovss.n1752 9.0005
R1803 iovss.n1824 iovss.n1752 9.0005
R1804 iovss.n1790 iovss.n1752 9.0005
R1805 iovss.n1827 iovss.n1752 9.0005
R1806 iovss.n1789 iovss.n1752 9.0005
R1807 iovss.n1830 iovss.n1752 9.0005
R1808 iovss.n1788 iovss.n1752 9.0005
R1809 iovss.n1832 iovss.n1752 9.0005
R1810 iovss.n1787 iovss.n1752 9.0005
R1811 iovss.n1835 iovss.n1752 9.0005
R1812 iovss.n1786 iovss.n1752 9.0005
R1813 iovss.n1837 iovss.n1752 9.0005
R1814 iovss.n1785 iovss.n1752 9.0005
R1815 iovss.n1840 iovss.n1752 9.0005
R1816 iovss.n1784 iovss.n1752 9.0005
R1817 iovss.n1841 iovss.n1752 9.0005
R1818 iovss.n1870 iovss.n1752 9.0005
R1819 iovss.n2290 iovss.n1752 9.0005
R1820 iovss.n2292 iovss.n1710 9.0005
R1821 iovss.n1801 iovss.n1710 9.0005
R1822 iovss.n1799 iovss.n1710 9.0005
R1823 iovss.n1804 iovss.n1710 9.0005
R1824 iovss.n1798 iovss.n1710 9.0005
R1825 iovss.n1807 iovss.n1710 9.0005
R1826 iovss.n1797 iovss.n1710 9.0005
R1827 iovss.n1809 iovss.n1710 9.0005
R1828 iovss.n1796 iovss.n1710 9.0005
R1829 iovss.n1812 iovss.n1710 9.0005
R1830 iovss.n1795 iovss.n1710 9.0005
R1831 iovss.n1814 iovss.n1710 9.0005
R1832 iovss.n1794 iovss.n1710 9.0005
R1833 iovss.n1817 iovss.n1710 9.0005
R1834 iovss.n1793 iovss.n1710 9.0005
R1835 iovss.n1819 iovss.n1710 9.0005
R1836 iovss.n1792 iovss.n1710 9.0005
R1837 iovss.n1822 iovss.n1710 9.0005
R1838 iovss.n1791 iovss.n1710 9.0005
R1839 iovss.n1824 iovss.n1710 9.0005
R1840 iovss.n1790 iovss.n1710 9.0005
R1841 iovss.n1827 iovss.n1710 9.0005
R1842 iovss.n1789 iovss.n1710 9.0005
R1843 iovss.n1830 iovss.n1710 9.0005
R1844 iovss.n1788 iovss.n1710 9.0005
R1845 iovss.n1832 iovss.n1710 9.0005
R1846 iovss.n1787 iovss.n1710 9.0005
R1847 iovss.n1835 iovss.n1710 9.0005
R1848 iovss.n1786 iovss.n1710 9.0005
R1849 iovss.n1837 iovss.n1710 9.0005
R1850 iovss.n1785 iovss.n1710 9.0005
R1851 iovss.n1840 iovss.n1710 9.0005
R1852 iovss.n1784 iovss.n1710 9.0005
R1853 iovss.n1841 iovss.n1710 9.0005
R1854 iovss.n1870 iovss.n1710 9.0005
R1855 iovss.n2290 iovss.n1710 9.0005
R1856 iovss.n2292 iovss.n1753 9.0005
R1857 iovss.n1801 iovss.n1753 9.0005
R1858 iovss.n1799 iovss.n1753 9.0005
R1859 iovss.n1804 iovss.n1753 9.0005
R1860 iovss.n1798 iovss.n1753 9.0005
R1861 iovss.n1807 iovss.n1753 9.0005
R1862 iovss.n1797 iovss.n1753 9.0005
R1863 iovss.n1809 iovss.n1753 9.0005
R1864 iovss.n1796 iovss.n1753 9.0005
R1865 iovss.n1812 iovss.n1753 9.0005
R1866 iovss.n1795 iovss.n1753 9.0005
R1867 iovss.n1814 iovss.n1753 9.0005
R1868 iovss.n1794 iovss.n1753 9.0005
R1869 iovss.n1817 iovss.n1753 9.0005
R1870 iovss.n1793 iovss.n1753 9.0005
R1871 iovss.n1819 iovss.n1753 9.0005
R1872 iovss.n1792 iovss.n1753 9.0005
R1873 iovss.n1822 iovss.n1753 9.0005
R1874 iovss.n1791 iovss.n1753 9.0005
R1875 iovss.n1824 iovss.n1753 9.0005
R1876 iovss.n1790 iovss.n1753 9.0005
R1877 iovss.n1827 iovss.n1753 9.0005
R1878 iovss.n1789 iovss.n1753 9.0005
R1879 iovss.n1830 iovss.n1753 9.0005
R1880 iovss.n1788 iovss.n1753 9.0005
R1881 iovss.n1832 iovss.n1753 9.0005
R1882 iovss.n1787 iovss.n1753 9.0005
R1883 iovss.n1835 iovss.n1753 9.0005
R1884 iovss.n1786 iovss.n1753 9.0005
R1885 iovss.n1837 iovss.n1753 9.0005
R1886 iovss.n1785 iovss.n1753 9.0005
R1887 iovss.n1840 iovss.n1753 9.0005
R1888 iovss.n1784 iovss.n1753 9.0005
R1889 iovss.n1841 iovss.n1753 9.0005
R1890 iovss.n1870 iovss.n1753 9.0005
R1891 iovss.n2290 iovss.n1753 9.0005
R1892 iovss.n2292 iovss.n1709 9.0005
R1893 iovss.n1801 iovss.n1709 9.0005
R1894 iovss.n1799 iovss.n1709 9.0005
R1895 iovss.n1804 iovss.n1709 9.0005
R1896 iovss.n1798 iovss.n1709 9.0005
R1897 iovss.n1807 iovss.n1709 9.0005
R1898 iovss.n1797 iovss.n1709 9.0005
R1899 iovss.n1809 iovss.n1709 9.0005
R1900 iovss.n1796 iovss.n1709 9.0005
R1901 iovss.n1812 iovss.n1709 9.0005
R1902 iovss.n1795 iovss.n1709 9.0005
R1903 iovss.n1814 iovss.n1709 9.0005
R1904 iovss.n1794 iovss.n1709 9.0005
R1905 iovss.n1817 iovss.n1709 9.0005
R1906 iovss.n1793 iovss.n1709 9.0005
R1907 iovss.n1819 iovss.n1709 9.0005
R1908 iovss.n1792 iovss.n1709 9.0005
R1909 iovss.n1822 iovss.n1709 9.0005
R1910 iovss.n1791 iovss.n1709 9.0005
R1911 iovss.n1824 iovss.n1709 9.0005
R1912 iovss.n1790 iovss.n1709 9.0005
R1913 iovss.n1827 iovss.n1709 9.0005
R1914 iovss.n1789 iovss.n1709 9.0005
R1915 iovss.n1830 iovss.n1709 9.0005
R1916 iovss.n1788 iovss.n1709 9.0005
R1917 iovss.n1832 iovss.n1709 9.0005
R1918 iovss.n1787 iovss.n1709 9.0005
R1919 iovss.n1835 iovss.n1709 9.0005
R1920 iovss.n1786 iovss.n1709 9.0005
R1921 iovss.n1837 iovss.n1709 9.0005
R1922 iovss.n1785 iovss.n1709 9.0005
R1923 iovss.n1840 iovss.n1709 9.0005
R1924 iovss.n1784 iovss.n1709 9.0005
R1925 iovss.n1841 iovss.n1709 9.0005
R1926 iovss.n1870 iovss.n1709 9.0005
R1927 iovss.n2290 iovss.n1709 9.0005
R1928 iovss.n2292 iovss.n1754 9.0005
R1929 iovss.n1801 iovss.n1754 9.0005
R1930 iovss.n1799 iovss.n1754 9.0005
R1931 iovss.n1804 iovss.n1754 9.0005
R1932 iovss.n1798 iovss.n1754 9.0005
R1933 iovss.n1807 iovss.n1754 9.0005
R1934 iovss.n1797 iovss.n1754 9.0005
R1935 iovss.n1809 iovss.n1754 9.0005
R1936 iovss.n1796 iovss.n1754 9.0005
R1937 iovss.n1812 iovss.n1754 9.0005
R1938 iovss.n1795 iovss.n1754 9.0005
R1939 iovss.n1814 iovss.n1754 9.0005
R1940 iovss.n1794 iovss.n1754 9.0005
R1941 iovss.n1817 iovss.n1754 9.0005
R1942 iovss.n1793 iovss.n1754 9.0005
R1943 iovss.n1819 iovss.n1754 9.0005
R1944 iovss.n1792 iovss.n1754 9.0005
R1945 iovss.n1822 iovss.n1754 9.0005
R1946 iovss.n1791 iovss.n1754 9.0005
R1947 iovss.n1824 iovss.n1754 9.0005
R1948 iovss.n1790 iovss.n1754 9.0005
R1949 iovss.n1827 iovss.n1754 9.0005
R1950 iovss.n1789 iovss.n1754 9.0005
R1951 iovss.n1830 iovss.n1754 9.0005
R1952 iovss.n1788 iovss.n1754 9.0005
R1953 iovss.n1832 iovss.n1754 9.0005
R1954 iovss.n1787 iovss.n1754 9.0005
R1955 iovss.n1835 iovss.n1754 9.0005
R1956 iovss.n1786 iovss.n1754 9.0005
R1957 iovss.n1837 iovss.n1754 9.0005
R1958 iovss.n1785 iovss.n1754 9.0005
R1959 iovss.n1840 iovss.n1754 9.0005
R1960 iovss.n1784 iovss.n1754 9.0005
R1961 iovss.n1841 iovss.n1754 9.0005
R1962 iovss.n1870 iovss.n1754 9.0005
R1963 iovss.n2290 iovss.n1754 9.0005
R1964 iovss.n2292 iovss.n1708 9.0005
R1965 iovss.n1801 iovss.n1708 9.0005
R1966 iovss.n1799 iovss.n1708 9.0005
R1967 iovss.n1804 iovss.n1708 9.0005
R1968 iovss.n1798 iovss.n1708 9.0005
R1969 iovss.n1807 iovss.n1708 9.0005
R1970 iovss.n1797 iovss.n1708 9.0005
R1971 iovss.n1809 iovss.n1708 9.0005
R1972 iovss.n1796 iovss.n1708 9.0005
R1973 iovss.n1812 iovss.n1708 9.0005
R1974 iovss.n1795 iovss.n1708 9.0005
R1975 iovss.n1814 iovss.n1708 9.0005
R1976 iovss.n1794 iovss.n1708 9.0005
R1977 iovss.n1817 iovss.n1708 9.0005
R1978 iovss.n1793 iovss.n1708 9.0005
R1979 iovss.n1819 iovss.n1708 9.0005
R1980 iovss.n1792 iovss.n1708 9.0005
R1981 iovss.n1822 iovss.n1708 9.0005
R1982 iovss.n1791 iovss.n1708 9.0005
R1983 iovss.n1824 iovss.n1708 9.0005
R1984 iovss.n1790 iovss.n1708 9.0005
R1985 iovss.n1827 iovss.n1708 9.0005
R1986 iovss.n1789 iovss.n1708 9.0005
R1987 iovss.n1830 iovss.n1708 9.0005
R1988 iovss.n1788 iovss.n1708 9.0005
R1989 iovss.n1832 iovss.n1708 9.0005
R1990 iovss.n1787 iovss.n1708 9.0005
R1991 iovss.n1835 iovss.n1708 9.0005
R1992 iovss.n1786 iovss.n1708 9.0005
R1993 iovss.n1837 iovss.n1708 9.0005
R1994 iovss.n1785 iovss.n1708 9.0005
R1995 iovss.n1840 iovss.n1708 9.0005
R1996 iovss.n1784 iovss.n1708 9.0005
R1997 iovss.n1841 iovss.n1708 9.0005
R1998 iovss.n1870 iovss.n1708 9.0005
R1999 iovss.n2290 iovss.n1708 9.0005
R2000 iovss.n2292 iovss.n1755 9.0005
R2001 iovss.n1801 iovss.n1755 9.0005
R2002 iovss.n1799 iovss.n1755 9.0005
R2003 iovss.n1804 iovss.n1755 9.0005
R2004 iovss.n1798 iovss.n1755 9.0005
R2005 iovss.n1807 iovss.n1755 9.0005
R2006 iovss.n1797 iovss.n1755 9.0005
R2007 iovss.n1809 iovss.n1755 9.0005
R2008 iovss.n1796 iovss.n1755 9.0005
R2009 iovss.n1812 iovss.n1755 9.0005
R2010 iovss.n1795 iovss.n1755 9.0005
R2011 iovss.n1814 iovss.n1755 9.0005
R2012 iovss.n1794 iovss.n1755 9.0005
R2013 iovss.n1817 iovss.n1755 9.0005
R2014 iovss.n1793 iovss.n1755 9.0005
R2015 iovss.n1819 iovss.n1755 9.0005
R2016 iovss.n1792 iovss.n1755 9.0005
R2017 iovss.n1822 iovss.n1755 9.0005
R2018 iovss.n1791 iovss.n1755 9.0005
R2019 iovss.n1824 iovss.n1755 9.0005
R2020 iovss.n1790 iovss.n1755 9.0005
R2021 iovss.n1827 iovss.n1755 9.0005
R2022 iovss.n1789 iovss.n1755 9.0005
R2023 iovss.n1830 iovss.n1755 9.0005
R2024 iovss.n1788 iovss.n1755 9.0005
R2025 iovss.n1832 iovss.n1755 9.0005
R2026 iovss.n1787 iovss.n1755 9.0005
R2027 iovss.n1835 iovss.n1755 9.0005
R2028 iovss.n1786 iovss.n1755 9.0005
R2029 iovss.n1837 iovss.n1755 9.0005
R2030 iovss.n1785 iovss.n1755 9.0005
R2031 iovss.n1840 iovss.n1755 9.0005
R2032 iovss.n1784 iovss.n1755 9.0005
R2033 iovss.n1841 iovss.n1755 9.0005
R2034 iovss.n1870 iovss.n1755 9.0005
R2035 iovss.n2290 iovss.n1755 9.0005
R2036 iovss.n2292 iovss.n1707 9.0005
R2037 iovss.n1801 iovss.n1707 9.0005
R2038 iovss.n1799 iovss.n1707 9.0005
R2039 iovss.n1804 iovss.n1707 9.0005
R2040 iovss.n1798 iovss.n1707 9.0005
R2041 iovss.n1807 iovss.n1707 9.0005
R2042 iovss.n1797 iovss.n1707 9.0005
R2043 iovss.n1809 iovss.n1707 9.0005
R2044 iovss.n1796 iovss.n1707 9.0005
R2045 iovss.n1812 iovss.n1707 9.0005
R2046 iovss.n1795 iovss.n1707 9.0005
R2047 iovss.n1814 iovss.n1707 9.0005
R2048 iovss.n1794 iovss.n1707 9.0005
R2049 iovss.n1817 iovss.n1707 9.0005
R2050 iovss.n1793 iovss.n1707 9.0005
R2051 iovss.n1819 iovss.n1707 9.0005
R2052 iovss.n1792 iovss.n1707 9.0005
R2053 iovss.n1822 iovss.n1707 9.0005
R2054 iovss.n1791 iovss.n1707 9.0005
R2055 iovss.n1824 iovss.n1707 9.0005
R2056 iovss.n1790 iovss.n1707 9.0005
R2057 iovss.n1827 iovss.n1707 9.0005
R2058 iovss.n1789 iovss.n1707 9.0005
R2059 iovss.n1830 iovss.n1707 9.0005
R2060 iovss.n1788 iovss.n1707 9.0005
R2061 iovss.n1832 iovss.n1707 9.0005
R2062 iovss.n1787 iovss.n1707 9.0005
R2063 iovss.n1835 iovss.n1707 9.0005
R2064 iovss.n1786 iovss.n1707 9.0005
R2065 iovss.n1837 iovss.n1707 9.0005
R2066 iovss.n1785 iovss.n1707 9.0005
R2067 iovss.n1840 iovss.n1707 9.0005
R2068 iovss.n1784 iovss.n1707 9.0005
R2069 iovss.n1841 iovss.n1707 9.0005
R2070 iovss.n1870 iovss.n1707 9.0005
R2071 iovss.n2290 iovss.n1707 9.0005
R2072 iovss.n2292 iovss.n1756 9.0005
R2073 iovss.n1801 iovss.n1756 9.0005
R2074 iovss.n1799 iovss.n1756 9.0005
R2075 iovss.n1804 iovss.n1756 9.0005
R2076 iovss.n1798 iovss.n1756 9.0005
R2077 iovss.n1807 iovss.n1756 9.0005
R2078 iovss.n1797 iovss.n1756 9.0005
R2079 iovss.n1809 iovss.n1756 9.0005
R2080 iovss.n1796 iovss.n1756 9.0005
R2081 iovss.n1812 iovss.n1756 9.0005
R2082 iovss.n1795 iovss.n1756 9.0005
R2083 iovss.n1814 iovss.n1756 9.0005
R2084 iovss.n1794 iovss.n1756 9.0005
R2085 iovss.n1817 iovss.n1756 9.0005
R2086 iovss.n1793 iovss.n1756 9.0005
R2087 iovss.n1819 iovss.n1756 9.0005
R2088 iovss.n1792 iovss.n1756 9.0005
R2089 iovss.n1822 iovss.n1756 9.0005
R2090 iovss.n1791 iovss.n1756 9.0005
R2091 iovss.n1824 iovss.n1756 9.0005
R2092 iovss.n1790 iovss.n1756 9.0005
R2093 iovss.n1827 iovss.n1756 9.0005
R2094 iovss.n1789 iovss.n1756 9.0005
R2095 iovss.n1830 iovss.n1756 9.0005
R2096 iovss.n1788 iovss.n1756 9.0005
R2097 iovss.n1832 iovss.n1756 9.0005
R2098 iovss.n1787 iovss.n1756 9.0005
R2099 iovss.n1835 iovss.n1756 9.0005
R2100 iovss.n1786 iovss.n1756 9.0005
R2101 iovss.n1837 iovss.n1756 9.0005
R2102 iovss.n1785 iovss.n1756 9.0005
R2103 iovss.n1840 iovss.n1756 9.0005
R2104 iovss.n1784 iovss.n1756 9.0005
R2105 iovss.n1841 iovss.n1756 9.0005
R2106 iovss.n1870 iovss.n1756 9.0005
R2107 iovss.n2290 iovss.n1756 9.0005
R2108 iovss.n2292 iovss.n1706 9.0005
R2109 iovss.n1801 iovss.n1706 9.0005
R2110 iovss.n1799 iovss.n1706 9.0005
R2111 iovss.n1804 iovss.n1706 9.0005
R2112 iovss.n1798 iovss.n1706 9.0005
R2113 iovss.n1807 iovss.n1706 9.0005
R2114 iovss.n1797 iovss.n1706 9.0005
R2115 iovss.n1809 iovss.n1706 9.0005
R2116 iovss.n1796 iovss.n1706 9.0005
R2117 iovss.n1812 iovss.n1706 9.0005
R2118 iovss.n1795 iovss.n1706 9.0005
R2119 iovss.n1814 iovss.n1706 9.0005
R2120 iovss.n1794 iovss.n1706 9.0005
R2121 iovss.n1817 iovss.n1706 9.0005
R2122 iovss.n1793 iovss.n1706 9.0005
R2123 iovss.n1819 iovss.n1706 9.0005
R2124 iovss.n1792 iovss.n1706 9.0005
R2125 iovss.n1822 iovss.n1706 9.0005
R2126 iovss.n1791 iovss.n1706 9.0005
R2127 iovss.n1824 iovss.n1706 9.0005
R2128 iovss.n1790 iovss.n1706 9.0005
R2129 iovss.n1827 iovss.n1706 9.0005
R2130 iovss.n1789 iovss.n1706 9.0005
R2131 iovss.n1830 iovss.n1706 9.0005
R2132 iovss.n1788 iovss.n1706 9.0005
R2133 iovss.n1832 iovss.n1706 9.0005
R2134 iovss.n1787 iovss.n1706 9.0005
R2135 iovss.n1835 iovss.n1706 9.0005
R2136 iovss.n1786 iovss.n1706 9.0005
R2137 iovss.n1837 iovss.n1706 9.0005
R2138 iovss.n1785 iovss.n1706 9.0005
R2139 iovss.n1840 iovss.n1706 9.0005
R2140 iovss.n1784 iovss.n1706 9.0005
R2141 iovss.n1841 iovss.n1706 9.0005
R2142 iovss.n1870 iovss.n1706 9.0005
R2143 iovss.n2290 iovss.n1706 9.0005
R2144 iovss.n2292 iovss.n2291 9.0005
R2145 iovss.n2291 iovss.n1801 9.0005
R2146 iovss.n2291 iovss.n1799 9.0005
R2147 iovss.n2291 iovss.n1804 9.0005
R2148 iovss.n2291 iovss.n1798 9.0005
R2149 iovss.n2291 iovss.n1807 9.0005
R2150 iovss.n2291 iovss.n1797 9.0005
R2151 iovss.n2291 iovss.n1809 9.0005
R2152 iovss.n2291 iovss.n1796 9.0005
R2153 iovss.n2291 iovss.n1812 9.0005
R2154 iovss.n2291 iovss.n1795 9.0005
R2155 iovss.n2291 iovss.n1814 9.0005
R2156 iovss.n2291 iovss.n1794 9.0005
R2157 iovss.n2291 iovss.n1817 9.0005
R2158 iovss.n2291 iovss.n1793 9.0005
R2159 iovss.n2291 iovss.n1819 9.0005
R2160 iovss.n2291 iovss.n1792 9.0005
R2161 iovss.n2291 iovss.n1822 9.0005
R2162 iovss.n2291 iovss.n1791 9.0005
R2163 iovss.n2291 iovss.n1824 9.0005
R2164 iovss.n2291 iovss.n1790 9.0005
R2165 iovss.n2291 iovss.n1827 9.0005
R2166 iovss.n2291 iovss.n1789 9.0005
R2167 iovss.n2291 iovss.n1830 9.0005
R2168 iovss.n2291 iovss.n1788 9.0005
R2169 iovss.n2291 iovss.n1832 9.0005
R2170 iovss.n2291 iovss.n1787 9.0005
R2171 iovss.n2291 iovss.n1835 9.0005
R2172 iovss.n2291 iovss.n1786 9.0005
R2173 iovss.n2291 iovss.n1837 9.0005
R2174 iovss.n2291 iovss.n1785 9.0005
R2175 iovss.n2291 iovss.n1840 9.0005
R2176 iovss.n2291 iovss.n1784 9.0005
R2177 iovss.n2291 iovss.n1841 9.0005
R2178 iovss.n2291 iovss.n1870 9.0005
R2179 iovss.n2291 iovss.n1783 9.0005
R2180 iovss.n2291 iovss.n2290 9.0005
R2181 iovss.n1961 iovss.n673 9.0005
R2182 iovss.n2121 iovss.n673 9.0005
R2183 iovss.n1949 iovss.n673 9.0005
R2184 iovss.n2126 iovss.n673 9.0005
R2185 iovss.n1947 iovss.n673 9.0005
R2186 iovss.n2131 iovss.n673 9.0005
R2187 iovss.n1945 iovss.n673 9.0005
R2188 iovss.n2162 iovss.n673 9.0005
R2189 iovss.n2241 iovss.n673 9.0005
R2190 iovss.n2243 iovss.n1918 9.0005
R2191 iovss.n1918 iovss.n1891 9.0005
R2192 iovss.n1958 iovss.n1918 9.0005
R2193 iovss.n2101 iovss.n1918 9.0005
R2194 iovss.n1956 iovss.n1918 9.0005
R2195 iovss.n2106 iovss.n1918 9.0005
R2196 iovss.n1954 iovss.n1918 9.0005
R2197 iovss.n2111 iovss.n1918 9.0005
R2198 iovss.n1952 iovss.n1918 9.0005
R2199 iovss.n2116 iovss.n1918 9.0005
R2200 iovss.n2162 iovss.n1918 9.0005
R2201 iovss.n2241 iovss.n1918 9.0005
R2202 iovss.n1961 iovss.n1916 9.0005
R2203 iovss.n2095 iovss.n1916 9.0005
R2204 iovss.n2243 iovss.n1916 9.0005
R2205 iovss.n1916 iovss.n1891 9.0005
R2206 iovss.n1960 iovss.n1916 9.0005
R2207 iovss.n2098 iovss.n1916 9.0005
R2208 iovss.n1958 iovss.n1916 9.0005
R2209 iovss.n2101 iovss.n1916 9.0005
R2210 iovss.n1957 iovss.n1916 9.0005
R2211 iovss.n2104 iovss.n1916 9.0005
R2212 iovss.n1956 iovss.n1916 9.0005
R2213 iovss.n2106 iovss.n1916 9.0005
R2214 iovss.n1955 iovss.n1916 9.0005
R2215 iovss.n2109 iovss.n1916 9.0005
R2216 iovss.n1954 iovss.n1916 9.0005
R2217 iovss.n2111 iovss.n1916 9.0005
R2218 iovss.n1953 iovss.n1916 9.0005
R2219 iovss.n2114 iovss.n1916 9.0005
R2220 iovss.n1952 iovss.n1916 9.0005
R2221 iovss.n2116 iovss.n1916 9.0005
R2222 iovss.n1951 iovss.n1916 9.0005
R2223 iovss.n2119 iovss.n1916 9.0005
R2224 iovss.n1950 iovss.n1916 9.0005
R2225 iovss.n2121 iovss.n1916 9.0005
R2226 iovss.n1949 iovss.n1916 9.0005
R2227 iovss.n2124 iovss.n1916 9.0005
R2228 iovss.n1948 iovss.n1916 9.0005
R2229 iovss.n2126 iovss.n1916 9.0005
R2230 iovss.n1947 iovss.n1916 9.0005
R2231 iovss.n2129 iovss.n1916 9.0005
R2232 iovss.n1946 iovss.n1916 9.0005
R2233 iovss.n2131 iovss.n1916 9.0005
R2234 iovss.n1945 iovss.n1916 9.0005
R2235 iovss.n2160 iovss.n1916 9.0005
R2236 iovss.n2162 iovss.n1916 9.0005
R2237 iovss.n2241 iovss.n1916 9.0005
R2238 iovss.n1961 iovss.n1919 9.0005
R2239 iovss.n2095 iovss.n1919 9.0005
R2240 iovss.n2243 iovss.n1919 9.0005
R2241 iovss.n1919 iovss.n1891 9.0005
R2242 iovss.n1960 iovss.n1919 9.0005
R2243 iovss.n2098 iovss.n1919 9.0005
R2244 iovss.n1958 iovss.n1919 9.0005
R2245 iovss.n2101 iovss.n1919 9.0005
R2246 iovss.n1957 iovss.n1919 9.0005
R2247 iovss.n2104 iovss.n1919 9.0005
R2248 iovss.n1956 iovss.n1919 9.0005
R2249 iovss.n2106 iovss.n1919 9.0005
R2250 iovss.n1955 iovss.n1919 9.0005
R2251 iovss.n2109 iovss.n1919 9.0005
R2252 iovss.n1954 iovss.n1919 9.0005
R2253 iovss.n2111 iovss.n1919 9.0005
R2254 iovss.n1953 iovss.n1919 9.0005
R2255 iovss.n2114 iovss.n1919 9.0005
R2256 iovss.n1952 iovss.n1919 9.0005
R2257 iovss.n2116 iovss.n1919 9.0005
R2258 iovss.n1951 iovss.n1919 9.0005
R2259 iovss.n2119 iovss.n1919 9.0005
R2260 iovss.n1950 iovss.n1919 9.0005
R2261 iovss.n2121 iovss.n1919 9.0005
R2262 iovss.n1949 iovss.n1919 9.0005
R2263 iovss.n2124 iovss.n1919 9.0005
R2264 iovss.n1948 iovss.n1919 9.0005
R2265 iovss.n2126 iovss.n1919 9.0005
R2266 iovss.n1947 iovss.n1919 9.0005
R2267 iovss.n2129 iovss.n1919 9.0005
R2268 iovss.n1946 iovss.n1919 9.0005
R2269 iovss.n2131 iovss.n1919 9.0005
R2270 iovss.n1945 iovss.n1919 9.0005
R2271 iovss.n2160 iovss.n1919 9.0005
R2272 iovss.n2162 iovss.n1919 9.0005
R2273 iovss.n2241 iovss.n1919 9.0005
R2274 iovss.n1961 iovss.n1915 9.0005
R2275 iovss.n2095 iovss.n1915 9.0005
R2276 iovss.n2243 iovss.n1915 9.0005
R2277 iovss.n1915 iovss.n1891 9.0005
R2278 iovss.n1960 iovss.n1915 9.0005
R2279 iovss.n2098 iovss.n1915 9.0005
R2280 iovss.n1958 iovss.n1915 9.0005
R2281 iovss.n2101 iovss.n1915 9.0005
R2282 iovss.n1957 iovss.n1915 9.0005
R2283 iovss.n2104 iovss.n1915 9.0005
R2284 iovss.n1956 iovss.n1915 9.0005
R2285 iovss.n2106 iovss.n1915 9.0005
R2286 iovss.n1955 iovss.n1915 9.0005
R2287 iovss.n2109 iovss.n1915 9.0005
R2288 iovss.n1954 iovss.n1915 9.0005
R2289 iovss.n2111 iovss.n1915 9.0005
R2290 iovss.n1953 iovss.n1915 9.0005
R2291 iovss.n2114 iovss.n1915 9.0005
R2292 iovss.n1952 iovss.n1915 9.0005
R2293 iovss.n2116 iovss.n1915 9.0005
R2294 iovss.n1951 iovss.n1915 9.0005
R2295 iovss.n2119 iovss.n1915 9.0005
R2296 iovss.n1950 iovss.n1915 9.0005
R2297 iovss.n2121 iovss.n1915 9.0005
R2298 iovss.n1949 iovss.n1915 9.0005
R2299 iovss.n2124 iovss.n1915 9.0005
R2300 iovss.n1948 iovss.n1915 9.0005
R2301 iovss.n2126 iovss.n1915 9.0005
R2302 iovss.n1947 iovss.n1915 9.0005
R2303 iovss.n2129 iovss.n1915 9.0005
R2304 iovss.n1946 iovss.n1915 9.0005
R2305 iovss.n2131 iovss.n1915 9.0005
R2306 iovss.n1945 iovss.n1915 9.0005
R2307 iovss.n2160 iovss.n1915 9.0005
R2308 iovss.n2162 iovss.n1915 9.0005
R2309 iovss.n2241 iovss.n1915 9.0005
R2310 iovss.n1961 iovss.n1920 9.0005
R2311 iovss.n2095 iovss.n1920 9.0005
R2312 iovss.n2243 iovss.n1920 9.0005
R2313 iovss.n1920 iovss.n1891 9.0005
R2314 iovss.n1960 iovss.n1920 9.0005
R2315 iovss.n2098 iovss.n1920 9.0005
R2316 iovss.n1958 iovss.n1920 9.0005
R2317 iovss.n2101 iovss.n1920 9.0005
R2318 iovss.n1957 iovss.n1920 9.0005
R2319 iovss.n2104 iovss.n1920 9.0005
R2320 iovss.n1956 iovss.n1920 9.0005
R2321 iovss.n2106 iovss.n1920 9.0005
R2322 iovss.n1955 iovss.n1920 9.0005
R2323 iovss.n2109 iovss.n1920 9.0005
R2324 iovss.n1954 iovss.n1920 9.0005
R2325 iovss.n2111 iovss.n1920 9.0005
R2326 iovss.n1953 iovss.n1920 9.0005
R2327 iovss.n2114 iovss.n1920 9.0005
R2328 iovss.n1952 iovss.n1920 9.0005
R2329 iovss.n2116 iovss.n1920 9.0005
R2330 iovss.n1951 iovss.n1920 9.0005
R2331 iovss.n2119 iovss.n1920 9.0005
R2332 iovss.n1950 iovss.n1920 9.0005
R2333 iovss.n2121 iovss.n1920 9.0005
R2334 iovss.n1949 iovss.n1920 9.0005
R2335 iovss.n2124 iovss.n1920 9.0005
R2336 iovss.n1948 iovss.n1920 9.0005
R2337 iovss.n2126 iovss.n1920 9.0005
R2338 iovss.n1947 iovss.n1920 9.0005
R2339 iovss.n2129 iovss.n1920 9.0005
R2340 iovss.n1946 iovss.n1920 9.0005
R2341 iovss.n2131 iovss.n1920 9.0005
R2342 iovss.n1945 iovss.n1920 9.0005
R2343 iovss.n2160 iovss.n1920 9.0005
R2344 iovss.n2162 iovss.n1920 9.0005
R2345 iovss.n2241 iovss.n1920 9.0005
R2346 iovss.n1961 iovss.n1914 9.0005
R2347 iovss.n2095 iovss.n1914 9.0005
R2348 iovss.n2243 iovss.n1914 9.0005
R2349 iovss.n1914 iovss.n1891 9.0005
R2350 iovss.n1960 iovss.n1914 9.0005
R2351 iovss.n2098 iovss.n1914 9.0005
R2352 iovss.n1958 iovss.n1914 9.0005
R2353 iovss.n2101 iovss.n1914 9.0005
R2354 iovss.n1957 iovss.n1914 9.0005
R2355 iovss.n2104 iovss.n1914 9.0005
R2356 iovss.n1956 iovss.n1914 9.0005
R2357 iovss.n2106 iovss.n1914 9.0005
R2358 iovss.n1955 iovss.n1914 9.0005
R2359 iovss.n2109 iovss.n1914 9.0005
R2360 iovss.n1954 iovss.n1914 9.0005
R2361 iovss.n2111 iovss.n1914 9.0005
R2362 iovss.n1953 iovss.n1914 9.0005
R2363 iovss.n2114 iovss.n1914 9.0005
R2364 iovss.n1952 iovss.n1914 9.0005
R2365 iovss.n2116 iovss.n1914 9.0005
R2366 iovss.n1951 iovss.n1914 9.0005
R2367 iovss.n2119 iovss.n1914 9.0005
R2368 iovss.n1950 iovss.n1914 9.0005
R2369 iovss.n2121 iovss.n1914 9.0005
R2370 iovss.n1949 iovss.n1914 9.0005
R2371 iovss.n2124 iovss.n1914 9.0005
R2372 iovss.n1948 iovss.n1914 9.0005
R2373 iovss.n2126 iovss.n1914 9.0005
R2374 iovss.n1947 iovss.n1914 9.0005
R2375 iovss.n2129 iovss.n1914 9.0005
R2376 iovss.n1946 iovss.n1914 9.0005
R2377 iovss.n2131 iovss.n1914 9.0005
R2378 iovss.n1945 iovss.n1914 9.0005
R2379 iovss.n2160 iovss.n1914 9.0005
R2380 iovss.n2162 iovss.n1914 9.0005
R2381 iovss.n2241 iovss.n1914 9.0005
R2382 iovss.n1961 iovss.n1921 9.0005
R2383 iovss.n2095 iovss.n1921 9.0005
R2384 iovss.n2243 iovss.n1921 9.0005
R2385 iovss.n1921 iovss.n1891 9.0005
R2386 iovss.n1960 iovss.n1921 9.0005
R2387 iovss.n2098 iovss.n1921 9.0005
R2388 iovss.n1958 iovss.n1921 9.0005
R2389 iovss.n2101 iovss.n1921 9.0005
R2390 iovss.n1957 iovss.n1921 9.0005
R2391 iovss.n2104 iovss.n1921 9.0005
R2392 iovss.n1956 iovss.n1921 9.0005
R2393 iovss.n2106 iovss.n1921 9.0005
R2394 iovss.n1955 iovss.n1921 9.0005
R2395 iovss.n2109 iovss.n1921 9.0005
R2396 iovss.n1954 iovss.n1921 9.0005
R2397 iovss.n2111 iovss.n1921 9.0005
R2398 iovss.n1953 iovss.n1921 9.0005
R2399 iovss.n2114 iovss.n1921 9.0005
R2400 iovss.n1952 iovss.n1921 9.0005
R2401 iovss.n2116 iovss.n1921 9.0005
R2402 iovss.n1951 iovss.n1921 9.0005
R2403 iovss.n2119 iovss.n1921 9.0005
R2404 iovss.n1950 iovss.n1921 9.0005
R2405 iovss.n2121 iovss.n1921 9.0005
R2406 iovss.n1949 iovss.n1921 9.0005
R2407 iovss.n2124 iovss.n1921 9.0005
R2408 iovss.n1948 iovss.n1921 9.0005
R2409 iovss.n2126 iovss.n1921 9.0005
R2410 iovss.n1947 iovss.n1921 9.0005
R2411 iovss.n2129 iovss.n1921 9.0005
R2412 iovss.n1946 iovss.n1921 9.0005
R2413 iovss.n2131 iovss.n1921 9.0005
R2414 iovss.n1945 iovss.n1921 9.0005
R2415 iovss.n2160 iovss.n1921 9.0005
R2416 iovss.n2162 iovss.n1921 9.0005
R2417 iovss.n2241 iovss.n1921 9.0005
R2418 iovss.n1961 iovss.n1913 9.0005
R2419 iovss.n2095 iovss.n1913 9.0005
R2420 iovss.n2243 iovss.n1913 9.0005
R2421 iovss.n1913 iovss.n1891 9.0005
R2422 iovss.n1960 iovss.n1913 9.0005
R2423 iovss.n2098 iovss.n1913 9.0005
R2424 iovss.n1958 iovss.n1913 9.0005
R2425 iovss.n2101 iovss.n1913 9.0005
R2426 iovss.n1957 iovss.n1913 9.0005
R2427 iovss.n2104 iovss.n1913 9.0005
R2428 iovss.n1956 iovss.n1913 9.0005
R2429 iovss.n2106 iovss.n1913 9.0005
R2430 iovss.n1955 iovss.n1913 9.0005
R2431 iovss.n2109 iovss.n1913 9.0005
R2432 iovss.n1954 iovss.n1913 9.0005
R2433 iovss.n2111 iovss.n1913 9.0005
R2434 iovss.n1953 iovss.n1913 9.0005
R2435 iovss.n2114 iovss.n1913 9.0005
R2436 iovss.n1952 iovss.n1913 9.0005
R2437 iovss.n2116 iovss.n1913 9.0005
R2438 iovss.n1951 iovss.n1913 9.0005
R2439 iovss.n2119 iovss.n1913 9.0005
R2440 iovss.n1950 iovss.n1913 9.0005
R2441 iovss.n2121 iovss.n1913 9.0005
R2442 iovss.n1949 iovss.n1913 9.0005
R2443 iovss.n2124 iovss.n1913 9.0005
R2444 iovss.n1948 iovss.n1913 9.0005
R2445 iovss.n2126 iovss.n1913 9.0005
R2446 iovss.n1947 iovss.n1913 9.0005
R2447 iovss.n2129 iovss.n1913 9.0005
R2448 iovss.n1946 iovss.n1913 9.0005
R2449 iovss.n2131 iovss.n1913 9.0005
R2450 iovss.n1945 iovss.n1913 9.0005
R2451 iovss.n2160 iovss.n1913 9.0005
R2452 iovss.n2162 iovss.n1913 9.0005
R2453 iovss.n2241 iovss.n1913 9.0005
R2454 iovss.n1961 iovss.n1922 9.0005
R2455 iovss.n2095 iovss.n1922 9.0005
R2456 iovss.n2243 iovss.n1922 9.0005
R2457 iovss.n1922 iovss.n1891 9.0005
R2458 iovss.n1960 iovss.n1922 9.0005
R2459 iovss.n2098 iovss.n1922 9.0005
R2460 iovss.n1958 iovss.n1922 9.0005
R2461 iovss.n2101 iovss.n1922 9.0005
R2462 iovss.n1957 iovss.n1922 9.0005
R2463 iovss.n2104 iovss.n1922 9.0005
R2464 iovss.n1956 iovss.n1922 9.0005
R2465 iovss.n2106 iovss.n1922 9.0005
R2466 iovss.n1955 iovss.n1922 9.0005
R2467 iovss.n2109 iovss.n1922 9.0005
R2468 iovss.n1954 iovss.n1922 9.0005
R2469 iovss.n2111 iovss.n1922 9.0005
R2470 iovss.n1953 iovss.n1922 9.0005
R2471 iovss.n2114 iovss.n1922 9.0005
R2472 iovss.n1952 iovss.n1922 9.0005
R2473 iovss.n2116 iovss.n1922 9.0005
R2474 iovss.n1951 iovss.n1922 9.0005
R2475 iovss.n2119 iovss.n1922 9.0005
R2476 iovss.n1950 iovss.n1922 9.0005
R2477 iovss.n2121 iovss.n1922 9.0005
R2478 iovss.n1949 iovss.n1922 9.0005
R2479 iovss.n2124 iovss.n1922 9.0005
R2480 iovss.n1948 iovss.n1922 9.0005
R2481 iovss.n2126 iovss.n1922 9.0005
R2482 iovss.n1947 iovss.n1922 9.0005
R2483 iovss.n2129 iovss.n1922 9.0005
R2484 iovss.n1946 iovss.n1922 9.0005
R2485 iovss.n2131 iovss.n1922 9.0005
R2486 iovss.n1945 iovss.n1922 9.0005
R2487 iovss.n2160 iovss.n1922 9.0005
R2488 iovss.n2162 iovss.n1922 9.0005
R2489 iovss.n2241 iovss.n1922 9.0005
R2490 iovss.n1961 iovss.n1912 9.0005
R2491 iovss.n2095 iovss.n1912 9.0005
R2492 iovss.n2243 iovss.n1912 9.0005
R2493 iovss.n1912 iovss.n1891 9.0005
R2494 iovss.n1960 iovss.n1912 9.0005
R2495 iovss.n2098 iovss.n1912 9.0005
R2496 iovss.n1958 iovss.n1912 9.0005
R2497 iovss.n2101 iovss.n1912 9.0005
R2498 iovss.n1957 iovss.n1912 9.0005
R2499 iovss.n2104 iovss.n1912 9.0005
R2500 iovss.n1956 iovss.n1912 9.0005
R2501 iovss.n2106 iovss.n1912 9.0005
R2502 iovss.n1955 iovss.n1912 9.0005
R2503 iovss.n2109 iovss.n1912 9.0005
R2504 iovss.n1954 iovss.n1912 9.0005
R2505 iovss.n2111 iovss.n1912 9.0005
R2506 iovss.n1953 iovss.n1912 9.0005
R2507 iovss.n2114 iovss.n1912 9.0005
R2508 iovss.n1952 iovss.n1912 9.0005
R2509 iovss.n2116 iovss.n1912 9.0005
R2510 iovss.n1951 iovss.n1912 9.0005
R2511 iovss.n2119 iovss.n1912 9.0005
R2512 iovss.n1950 iovss.n1912 9.0005
R2513 iovss.n2121 iovss.n1912 9.0005
R2514 iovss.n1949 iovss.n1912 9.0005
R2515 iovss.n2124 iovss.n1912 9.0005
R2516 iovss.n1948 iovss.n1912 9.0005
R2517 iovss.n2126 iovss.n1912 9.0005
R2518 iovss.n1947 iovss.n1912 9.0005
R2519 iovss.n2129 iovss.n1912 9.0005
R2520 iovss.n1946 iovss.n1912 9.0005
R2521 iovss.n2131 iovss.n1912 9.0005
R2522 iovss.n1945 iovss.n1912 9.0005
R2523 iovss.n2160 iovss.n1912 9.0005
R2524 iovss.n2162 iovss.n1912 9.0005
R2525 iovss.n2241 iovss.n1912 9.0005
R2526 iovss.n1961 iovss.n1923 9.0005
R2527 iovss.n2095 iovss.n1923 9.0005
R2528 iovss.n2243 iovss.n1923 9.0005
R2529 iovss.n1923 iovss.n1891 9.0005
R2530 iovss.n1960 iovss.n1923 9.0005
R2531 iovss.n2098 iovss.n1923 9.0005
R2532 iovss.n1958 iovss.n1923 9.0005
R2533 iovss.n2101 iovss.n1923 9.0005
R2534 iovss.n1957 iovss.n1923 9.0005
R2535 iovss.n2104 iovss.n1923 9.0005
R2536 iovss.n1956 iovss.n1923 9.0005
R2537 iovss.n2106 iovss.n1923 9.0005
R2538 iovss.n1955 iovss.n1923 9.0005
R2539 iovss.n2109 iovss.n1923 9.0005
R2540 iovss.n1954 iovss.n1923 9.0005
R2541 iovss.n2111 iovss.n1923 9.0005
R2542 iovss.n1953 iovss.n1923 9.0005
R2543 iovss.n2114 iovss.n1923 9.0005
R2544 iovss.n1952 iovss.n1923 9.0005
R2545 iovss.n2116 iovss.n1923 9.0005
R2546 iovss.n1951 iovss.n1923 9.0005
R2547 iovss.n2119 iovss.n1923 9.0005
R2548 iovss.n1950 iovss.n1923 9.0005
R2549 iovss.n2121 iovss.n1923 9.0005
R2550 iovss.n1949 iovss.n1923 9.0005
R2551 iovss.n2124 iovss.n1923 9.0005
R2552 iovss.n1948 iovss.n1923 9.0005
R2553 iovss.n2126 iovss.n1923 9.0005
R2554 iovss.n1947 iovss.n1923 9.0005
R2555 iovss.n2129 iovss.n1923 9.0005
R2556 iovss.n1946 iovss.n1923 9.0005
R2557 iovss.n2131 iovss.n1923 9.0005
R2558 iovss.n1945 iovss.n1923 9.0005
R2559 iovss.n2160 iovss.n1923 9.0005
R2560 iovss.n2162 iovss.n1923 9.0005
R2561 iovss.n2241 iovss.n1923 9.0005
R2562 iovss.n1961 iovss.n1911 9.0005
R2563 iovss.n2095 iovss.n1911 9.0005
R2564 iovss.n2243 iovss.n1911 9.0005
R2565 iovss.n1911 iovss.n1891 9.0005
R2566 iovss.n1960 iovss.n1911 9.0005
R2567 iovss.n2098 iovss.n1911 9.0005
R2568 iovss.n1958 iovss.n1911 9.0005
R2569 iovss.n2101 iovss.n1911 9.0005
R2570 iovss.n1957 iovss.n1911 9.0005
R2571 iovss.n2104 iovss.n1911 9.0005
R2572 iovss.n1956 iovss.n1911 9.0005
R2573 iovss.n2106 iovss.n1911 9.0005
R2574 iovss.n1955 iovss.n1911 9.0005
R2575 iovss.n2109 iovss.n1911 9.0005
R2576 iovss.n1954 iovss.n1911 9.0005
R2577 iovss.n2111 iovss.n1911 9.0005
R2578 iovss.n1953 iovss.n1911 9.0005
R2579 iovss.n2114 iovss.n1911 9.0005
R2580 iovss.n1952 iovss.n1911 9.0005
R2581 iovss.n2116 iovss.n1911 9.0005
R2582 iovss.n1951 iovss.n1911 9.0005
R2583 iovss.n2119 iovss.n1911 9.0005
R2584 iovss.n1950 iovss.n1911 9.0005
R2585 iovss.n2121 iovss.n1911 9.0005
R2586 iovss.n1949 iovss.n1911 9.0005
R2587 iovss.n2124 iovss.n1911 9.0005
R2588 iovss.n1948 iovss.n1911 9.0005
R2589 iovss.n2126 iovss.n1911 9.0005
R2590 iovss.n1947 iovss.n1911 9.0005
R2591 iovss.n2129 iovss.n1911 9.0005
R2592 iovss.n1946 iovss.n1911 9.0005
R2593 iovss.n2131 iovss.n1911 9.0005
R2594 iovss.n1945 iovss.n1911 9.0005
R2595 iovss.n2160 iovss.n1911 9.0005
R2596 iovss.n2162 iovss.n1911 9.0005
R2597 iovss.n2241 iovss.n1911 9.0005
R2598 iovss.n1961 iovss.n1924 9.0005
R2599 iovss.n2095 iovss.n1924 9.0005
R2600 iovss.n2243 iovss.n1924 9.0005
R2601 iovss.n1924 iovss.n1891 9.0005
R2602 iovss.n1960 iovss.n1924 9.0005
R2603 iovss.n2098 iovss.n1924 9.0005
R2604 iovss.n1958 iovss.n1924 9.0005
R2605 iovss.n2101 iovss.n1924 9.0005
R2606 iovss.n1957 iovss.n1924 9.0005
R2607 iovss.n2104 iovss.n1924 9.0005
R2608 iovss.n1956 iovss.n1924 9.0005
R2609 iovss.n2106 iovss.n1924 9.0005
R2610 iovss.n1955 iovss.n1924 9.0005
R2611 iovss.n2109 iovss.n1924 9.0005
R2612 iovss.n1954 iovss.n1924 9.0005
R2613 iovss.n2111 iovss.n1924 9.0005
R2614 iovss.n1953 iovss.n1924 9.0005
R2615 iovss.n2114 iovss.n1924 9.0005
R2616 iovss.n1952 iovss.n1924 9.0005
R2617 iovss.n2116 iovss.n1924 9.0005
R2618 iovss.n1951 iovss.n1924 9.0005
R2619 iovss.n2119 iovss.n1924 9.0005
R2620 iovss.n1950 iovss.n1924 9.0005
R2621 iovss.n2121 iovss.n1924 9.0005
R2622 iovss.n1949 iovss.n1924 9.0005
R2623 iovss.n2124 iovss.n1924 9.0005
R2624 iovss.n1948 iovss.n1924 9.0005
R2625 iovss.n2126 iovss.n1924 9.0005
R2626 iovss.n1947 iovss.n1924 9.0005
R2627 iovss.n2129 iovss.n1924 9.0005
R2628 iovss.n1946 iovss.n1924 9.0005
R2629 iovss.n2131 iovss.n1924 9.0005
R2630 iovss.n1945 iovss.n1924 9.0005
R2631 iovss.n2160 iovss.n1924 9.0005
R2632 iovss.n2162 iovss.n1924 9.0005
R2633 iovss.n2241 iovss.n1924 9.0005
R2634 iovss.n1961 iovss.n1910 9.0005
R2635 iovss.n2095 iovss.n1910 9.0005
R2636 iovss.n2243 iovss.n1910 9.0005
R2637 iovss.n1910 iovss.n1891 9.0005
R2638 iovss.n1960 iovss.n1910 9.0005
R2639 iovss.n2098 iovss.n1910 9.0005
R2640 iovss.n1958 iovss.n1910 9.0005
R2641 iovss.n2101 iovss.n1910 9.0005
R2642 iovss.n1957 iovss.n1910 9.0005
R2643 iovss.n2104 iovss.n1910 9.0005
R2644 iovss.n1956 iovss.n1910 9.0005
R2645 iovss.n2106 iovss.n1910 9.0005
R2646 iovss.n1955 iovss.n1910 9.0005
R2647 iovss.n2109 iovss.n1910 9.0005
R2648 iovss.n1954 iovss.n1910 9.0005
R2649 iovss.n2111 iovss.n1910 9.0005
R2650 iovss.n1953 iovss.n1910 9.0005
R2651 iovss.n2114 iovss.n1910 9.0005
R2652 iovss.n1952 iovss.n1910 9.0005
R2653 iovss.n2116 iovss.n1910 9.0005
R2654 iovss.n1951 iovss.n1910 9.0005
R2655 iovss.n2119 iovss.n1910 9.0005
R2656 iovss.n1950 iovss.n1910 9.0005
R2657 iovss.n2121 iovss.n1910 9.0005
R2658 iovss.n1949 iovss.n1910 9.0005
R2659 iovss.n2124 iovss.n1910 9.0005
R2660 iovss.n1948 iovss.n1910 9.0005
R2661 iovss.n2126 iovss.n1910 9.0005
R2662 iovss.n1947 iovss.n1910 9.0005
R2663 iovss.n2129 iovss.n1910 9.0005
R2664 iovss.n1946 iovss.n1910 9.0005
R2665 iovss.n2131 iovss.n1910 9.0005
R2666 iovss.n1945 iovss.n1910 9.0005
R2667 iovss.n2160 iovss.n1910 9.0005
R2668 iovss.n2162 iovss.n1910 9.0005
R2669 iovss.n2241 iovss.n1910 9.0005
R2670 iovss.n1961 iovss.n1925 9.0005
R2671 iovss.n2095 iovss.n1925 9.0005
R2672 iovss.n2243 iovss.n1925 9.0005
R2673 iovss.n1925 iovss.n1891 9.0005
R2674 iovss.n1960 iovss.n1925 9.0005
R2675 iovss.n2098 iovss.n1925 9.0005
R2676 iovss.n1958 iovss.n1925 9.0005
R2677 iovss.n2101 iovss.n1925 9.0005
R2678 iovss.n1957 iovss.n1925 9.0005
R2679 iovss.n2104 iovss.n1925 9.0005
R2680 iovss.n1956 iovss.n1925 9.0005
R2681 iovss.n2106 iovss.n1925 9.0005
R2682 iovss.n1955 iovss.n1925 9.0005
R2683 iovss.n2109 iovss.n1925 9.0005
R2684 iovss.n1954 iovss.n1925 9.0005
R2685 iovss.n2111 iovss.n1925 9.0005
R2686 iovss.n1953 iovss.n1925 9.0005
R2687 iovss.n2114 iovss.n1925 9.0005
R2688 iovss.n1952 iovss.n1925 9.0005
R2689 iovss.n2116 iovss.n1925 9.0005
R2690 iovss.n1951 iovss.n1925 9.0005
R2691 iovss.n2119 iovss.n1925 9.0005
R2692 iovss.n1950 iovss.n1925 9.0005
R2693 iovss.n2121 iovss.n1925 9.0005
R2694 iovss.n1949 iovss.n1925 9.0005
R2695 iovss.n2124 iovss.n1925 9.0005
R2696 iovss.n1948 iovss.n1925 9.0005
R2697 iovss.n2126 iovss.n1925 9.0005
R2698 iovss.n1947 iovss.n1925 9.0005
R2699 iovss.n2129 iovss.n1925 9.0005
R2700 iovss.n1946 iovss.n1925 9.0005
R2701 iovss.n2131 iovss.n1925 9.0005
R2702 iovss.n1945 iovss.n1925 9.0005
R2703 iovss.n2160 iovss.n1925 9.0005
R2704 iovss.n2162 iovss.n1925 9.0005
R2705 iovss.n2241 iovss.n1925 9.0005
R2706 iovss.n1961 iovss.n1909 9.0005
R2707 iovss.n2095 iovss.n1909 9.0005
R2708 iovss.n2243 iovss.n1909 9.0005
R2709 iovss.n1909 iovss.n1891 9.0005
R2710 iovss.n1960 iovss.n1909 9.0005
R2711 iovss.n2098 iovss.n1909 9.0005
R2712 iovss.n1958 iovss.n1909 9.0005
R2713 iovss.n2101 iovss.n1909 9.0005
R2714 iovss.n1957 iovss.n1909 9.0005
R2715 iovss.n2104 iovss.n1909 9.0005
R2716 iovss.n1956 iovss.n1909 9.0005
R2717 iovss.n2106 iovss.n1909 9.0005
R2718 iovss.n1955 iovss.n1909 9.0005
R2719 iovss.n2109 iovss.n1909 9.0005
R2720 iovss.n1954 iovss.n1909 9.0005
R2721 iovss.n2111 iovss.n1909 9.0005
R2722 iovss.n1953 iovss.n1909 9.0005
R2723 iovss.n2114 iovss.n1909 9.0005
R2724 iovss.n1952 iovss.n1909 9.0005
R2725 iovss.n2116 iovss.n1909 9.0005
R2726 iovss.n1951 iovss.n1909 9.0005
R2727 iovss.n2119 iovss.n1909 9.0005
R2728 iovss.n1950 iovss.n1909 9.0005
R2729 iovss.n2121 iovss.n1909 9.0005
R2730 iovss.n1949 iovss.n1909 9.0005
R2731 iovss.n2124 iovss.n1909 9.0005
R2732 iovss.n1948 iovss.n1909 9.0005
R2733 iovss.n2126 iovss.n1909 9.0005
R2734 iovss.n1947 iovss.n1909 9.0005
R2735 iovss.n2129 iovss.n1909 9.0005
R2736 iovss.n1946 iovss.n1909 9.0005
R2737 iovss.n2131 iovss.n1909 9.0005
R2738 iovss.n1945 iovss.n1909 9.0005
R2739 iovss.n2160 iovss.n1909 9.0005
R2740 iovss.n2162 iovss.n1909 9.0005
R2741 iovss.n2241 iovss.n1909 9.0005
R2742 iovss.n1961 iovss.n1926 9.0005
R2743 iovss.n2095 iovss.n1926 9.0005
R2744 iovss.n2243 iovss.n1926 9.0005
R2745 iovss.n1926 iovss.n1891 9.0005
R2746 iovss.n1960 iovss.n1926 9.0005
R2747 iovss.n2098 iovss.n1926 9.0005
R2748 iovss.n1958 iovss.n1926 9.0005
R2749 iovss.n2101 iovss.n1926 9.0005
R2750 iovss.n1957 iovss.n1926 9.0005
R2751 iovss.n2104 iovss.n1926 9.0005
R2752 iovss.n1956 iovss.n1926 9.0005
R2753 iovss.n2106 iovss.n1926 9.0005
R2754 iovss.n1955 iovss.n1926 9.0005
R2755 iovss.n2109 iovss.n1926 9.0005
R2756 iovss.n1954 iovss.n1926 9.0005
R2757 iovss.n2111 iovss.n1926 9.0005
R2758 iovss.n1953 iovss.n1926 9.0005
R2759 iovss.n2114 iovss.n1926 9.0005
R2760 iovss.n1952 iovss.n1926 9.0005
R2761 iovss.n2116 iovss.n1926 9.0005
R2762 iovss.n1951 iovss.n1926 9.0005
R2763 iovss.n2119 iovss.n1926 9.0005
R2764 iovss.n1950 iovss.n1926 9.0005
R2765 iovss.n2121 iovss.n1926 9.0005
R2766 iovss.n1949 iovss.n1926 9.0005
R2767 iovss.n2124 iovss.n1926 9.0005
R2768 iovss.n1948 iovss.n1926 9.0005
R2769 iovss.n2126 iovss.n1926 9.0005
R2770 iovss.n1947 iovss.n1926 9.0005
R2771 iovss.n2129 iovss.n1926 9.0005
R2772 iovss.n1946 iovss.n1926 9.0005
R2773 iovss.n2131 iovss.n1926 9.0005
R2774 iovss.n1945 iovss.n1926 9.0005
R2775 iovss.n2160 iovss.n1926 9.0005
R2776 iovss.n2162 iovss.n1926 9.0005
R2777 iovss.n2241 iovss.n1926 9.0005
R2778 iovss.n1961 iovss.n1908 9.0005
R2779 iovss.n2095 iovss.n1908 9.0005
R2780 iovss.n2243 iovss.n1908 9.0005
R2781 iovss.n1908 iovss.n1891 9.0005
R2782 iovss.n1960 iovss.n1908 9.0005
R2783 iovss.n2098 iovss.n1908 9.0005
R2784 iovss.n1958 iovss.n1908 9.0005
R2785 iovss.n2101 iovss.n1908 9.0005
R2786 iovss.n1957 iovss.n1908 9.0005
R2787 iovss.n2104 iovss.n1908 9.0005
R2788 iovss.n1956 iovss.n1908 9.0005
R2789 iovss.n2106 iovss.n1908 9.0005
R2790 iovss.n1955 iovss.n1908 9.0005
R2791 iovss.n2109 iovss.n1908 9.0005
R2792 iovss.n1954 iovss.n1908 9.0005
R2793 iovss.n2111 iovss.n1908 9.0005
R2794 iovss.n1953 iovss.n1908 9.0005
R2795 iovss.n2114 iovss.n1908 9.0005
R2796 iovss.n1952 iovss.n1908 9.0005
R2797 iovss.n2116 iovss.n1908 9.0005
R2798 iovss.n1951 iovss.n1908 9.0005
R2799 iovss.n2119 iovss.n1908 9.0005
R2800 iovss.n1950 iovss.n1908 9.0005
R2801 iovss.n2121 iovss.n1908 9.0005
R2802 iovss.n1949 iovss.n1908 9.0005
R2803 iovss.n2124 iovss.n1908 9.0005
R2804 iovss.n1948 iovss.n1908 9.0005
R2805 iovss.n2126 iovss.n1908 9.0005
R2806 iovss.n1947 iovss.n1908 9.0005
R2807 iovss.n2129 iovss.n1908 9.0005
R2808 iovss.n1946 iovss.n1908 9.0005
R2809 iovss.n2131 iovss.n1908 9.0005
R2810 iovss.n1945 iovss.n1908 9.0005
R2811 iovss.n2160 iovss.n1908 9.0005
R2812 iovss.n2162 iovss.n1908 9.0005
R2813 iovss.n2241 iovss.n1908 9.0005
R2814 iovss.n1961 iovss.n1927 9.0005
R2815 iovss.n2095 iovss.n1927 9.0005
R2816 iovss.n2243 iovss.n1927 9.0005
R2817 iovss.n1927 iovss.n1891 9.0005
R2818 iovss.n1960 iovss.n1927 9.0005
R2819 iovss.n2098 iovss.n1927 9.0005
R2820 iovss.n1958 iovss.n1927 9.0005
R2821 iovss.n2101 iovss.n1927 9.0005
R2822 iovss.n1957 iovss.n1927 9.0005
R2823 iovss.n2104 iovss.n1927 9.0005
R2824 iovss.n1956 iovss.n1927 9.0005
R2825 iovss.n2106 iovss.n1927 9.0005
R2826 iovss.n1955 iovss.n1927 9.0005
R2827 iovss.n2109 iovss.n1927 9.0005
R2828 iovss.n1954 iovss.n1927 9.0005
R2829 iovss.n2111 iovss.n1927 9.0005
R2830 iovss.n1953 iovss.n1927 9.0005
R2831 iovss.n2114 iovss.n1927 9.0005
R2832 iovss.n1952 iovss.n1927 9.0005
R2833 iovss.n2116 iovss.n1927 9.0005
R2834 iovss.n1951 iovss.n1927 9.0005
R2835 iovss.n2119 iovss.n1927 9.0005
R2836 iovss.n1950 iovss.n1927 9.0005
R2837 iovss.n2121 iovss.n1927 9.0005
R2838 iovss.n1949 iovss.n1927 9.0005
R2839 iovss.n2124 iovss.n1927 9.0005
R2840 iovss.n1948 iovss.n1927 9.0005
R2841 iovss.n2126 iovss.n1927 9.0005
R2842 iovss.n1947 iovss.n1927 9.0005
R2843 iovss.n2129 iovss.n1927 9.0005
R2844 iovss.n1946 iovss.n1927 9.0005
R2845 iovss.n2131 iovss.n1927 9.0005
R2846 iovss.n1945 iovss.n1927 9.0005
R2847 iovss.n2160 iovss.n1927 9.0005
R2848 iovss.n2162 iovss.n1927 9.0005
R2849 iovss.n2241 iovss.n1927 9.0005
R2850 iovss.n1961 iovss.n1907 9.0005
R2851 iovss.n2095 iovss.n1907 9.0005
R2852 iovss.n2243 iovss.n1907 9.0005
R2853 iovss.n1907 iovss.n1891 9.0005
R2854 iovss.n1960 iovss.n1907 9.0005
R2855 iovss.n2098 iovss.n1907 9.0005
R2856 iovss.n1958 iovss.n1907 9.0005
R2857 iovss.n2101 iovss.n1907 9.0005
R2858 iovss.n1957 iovss.n1907 9.0005
R2859 iovss.n2104 iovss.n1907 9.0005
R2860 iovss.n1956 iovss.n1907 9.0005
R2861 iovss.n2106 iovss.n1907 9.0005
R2862 iovss.n1955 iovss.n1907 9.0005
R2863 iovss.n2109 iovss.n1907 9.0005
R2864 iovss.n1954 iovss.n1907 9.0005
R2865 iovss.n2111 iovss.n1907 9.0005
R2866 iovss.n1953 iovss.n1907 9.0005
R2867 iovss.n2114 iovss.n1907 9.0005
R2868 iovss.n1952 iovss.n1907 9.0005
R2869 iovss.n2116 iovss.n1907 9.0005
R2870 iovss.n1951 iovss.n1907 9.0005
R2871 iovss.n2119 iovss.n1907 9.0005
R2872 iovss.n1950 iovss.n1907 9.0005
R2873 iovss.n2121 iovss.n1907 9.0005
R2874 iovss.n1949 iovss.n1907 9.0005
R2875 iovss.n2124 iovss.n1907 9.0005
R2876 iovss.n1948 iovss.n1907 9.0005
R2877 iovss.n2126 iovss.n1907 9.0005
R2878 iovss.n1947 iovss.n1907 9.0005
R2879 iovss.n2129 iovss.n1907 9.0005
R2880 iovss.n1946 iovss.n1907 9.0005
R2881 iovss.n2131 iovss.n1907 9.0005
R2882 iovss.n1945 iovss.n1907 9.0005
R2883 iovss.n2160 iovss.n1907 9.0005
R2884 iovss.n2162 iovss.n1907 9.0005
R2885 iovss.n2241 iovss.n1907 9.0005
R2886 iovss.n1961 iovss.n1928 9.0005
R2887 iovss.n2095 iovss.n1928 9.0005
R2888 iovss.n2243 iovss.n1928 9.0005
R2889 iovss.n1928 iovss.n1891 9.0005
R2890 iovss.n1960 iovss.n1928 9.0005
R2891 iovss.n2098 iovss.n1928 9.0005
R2892 iovss.n1958 iovss.n1928 9.0005
R2893 iovss.n2101 iovss.n1928 9.0005
R2894 iovss.n1957 iovss.n1928 9.0005
R2895 iovss.n2104 iovss.n1928 9.0005
R2896 iovss.n1956 iovss.n1928 9.0005
R2897 iovss.n2106 iovss.n1928 9.0005
R2898 iovss.n1955 iovss.n1928 9.0005
R2899 iovss.n2109 iovss.n1928 9.0005
R2900 iovss.n1954 iovss.n1928 9.0005
R2901 iovss.n2111 iovss.n1928 9.0005
R2902 iovss.n1953 iovss.n1928 9.0005
R2903 iovss.n2114 iovss.n1928 9.0005
R2904 iovss.n1952 iovss.n1928 9.0005
R2905 iovss.n2116 iovss.n1928 9.0005
R2906 iovss.n1951 iovss.n1928 9.0005
R2907 iovss.n2119 iovss.n1928 9.0005
R2908 iovss.n1950 iovss.n1928 9.0005
R2909 iovss.n2121 iovss.n1928 9.0005
R2910 iovss.n1949 iovss.n1928 9.0005
R2911 iovss.n2124 iovss.n1928 9.0005
R2912 iovss.n1948 iovss.n1928 9.0005
R2913 iovss.n2126 iovss.n1928 9.0005
R2914 iovss.n1947 iovss.n1928 9.0005
R2915 iovss.n2129 iovss.n1928 9.0005
R2916 iovss.n1946 iovss.n1928 9.0005
R2917 iovss.n2131 iovss.n1928 9.0005
R2918 iovss.n1945 iovss.n1928 9.0005
R2919 iovss.n2160 iovss.n1928 9.0005
R2920 iovss.n2162 iovss.n1928 9.0005
R2921 iovss.n2241 iovss.n1928 9.0005
R2922 iovss.n1961 iovss.n1906 9.0005
R2923 iovss.n2095 iovss.n1906 9.0005
R2924 iovss.n2243 iovss.n1906 9.0005
R2925 iovss.n1906 iovss.n1891 9.0005
R2926 iovss.n1960 iovss.n1906 9.0005
R2927 iovss.n2098 iovss.n1906 9.0005
R2928 iovss.n1958 iovss.n1906 9.0005
R2929 iovss.n2101 iovss.n1906 9.0005
R2930 iovss.n1957 iovss.n1906 9.0005
R2931 iovss.n2104 iovss.n1906 9.0005
R2932 iovss.n1956 iovss.n1906 9.0005
R2933 iovss.n2106 iovss.n1906 9.0005
R2934 iovss.n1955 iovss.n1906 9.0005
R2935 iovss.n2109 iovss.n1906 9.0005
R2936 iovss.n1954 iovss.n1906 9.0005
R2937 iovss.n2111 iovss.n1906 9.0005
R2938 iovss.n1953 iovss.n1906 9.0005
R2939 iovss.n2114 iovss.n1906 9.0005
R2940 iovss.n1952 iovss.n1906 9.0005
R2941 iovss.n2116 iovss.n1906 9.0005
R2942 iovss.n1951 iovss.n1906 9.0005
R2943 iovss.n2119 iovss.n1906 9.0005
R2944 iovss.n1950 iovss.n1906 9.0005
R2945 iovss.n2121 iovss.n1906 9.0005
R2946 iovss.n1949 iovss.n1906 9.0005
R2947 iovss.n2124 iovss.n1906 9.0005
R2948 iovss.n1948 iovss.n1906 9.0005
R2949 iovss.n2126 iovss.n1906 9.0005
R2950 iovss.n1947 iovss.n1906 9.0005
R2951 iovss.n2129 iovss.n1906 9.0005
R2952 iovss.n1946 iovss.n1906 9.0005
R2953 iovss.n2131 iovss.n1906 9.0005
R2954 iovss.n1945 iovss.n1906 9.0005
R2955 iovss.n2160 iovss.n1906 9.0005
R2956 iovss.n2162 iovss.n1906 9.0005
R2957 iovss.n2241 iovss.n1906 9.0005
R2958 iovss.n1961 iovss.n1929 9.0005
R2959 iovss.n2095 iovss.n1929 9.0005
R2960 iovss.n2243 iovss.n1929 9.0005
R2961 iovss.n1929 iovss.n1891 9.0005
R2962 iovss.n1960 iovss.n1929 9.0005
R2963 iovss.n2098 iovss.n1929 9.0005
R2964 iovss.n1958 iovss.n1929 9.0005
R2965 iovss.n2101 iovss.n1929 9.0005
R2966 iovss.n1957 iovss.n1929 9.0005
R2967 iovss.n2104 iovss.n1929 9.0005
R2968 iovss.n1956 iovss.n1929 9.0005
R2969 iovss.n2106 iovss.n1929 9.0005
R2970 iovss.n1955 iovss.n1929 9.0005
R2971 iovss.n2109 iovss.n1929 9.0005
R2972 iovss.n1954 iovss.n1929 9.0005
R2973 iovss.n2111 iovss.n1929 9.0005
R2974 iovss.n1953 iovss.n1929 9.0005
R2975 iovss.n2114 iovss.n1929 9.0005
R2976 iovss.n1952 iovss.n1929 9.0005
R2977 iovss.n2116 iovss.n1929 9.0005
R2978 iovss.n1951 iovss.n1929 9.0005
R2979 iovss.n2119 iovss.n1929 9.0005
R2980 iovss.n1950 iovss.n1929 9.0005
R2981 iovss.n2121 iovss.n1929 9.0005
R2982 iovss.n1949 iovss.n1929 9.0005
R2983 iovss.n2124 iovss.n1929 9.0005
R2984 iovss.n1948 iovss.n1929 9.0005
R2985 iovss.n2126 iovss.n1929 9.0005
R2986 iovss.n1947 iovss.n1929 9.0005
R2987 iovss.n2129 iovss.n1929 9.0005
R2988 iovss.n1946 iovss.n1929 9.0005
R2989 iovss.n2131 iovss.n1929 9.0005
R2990 iovss.n1945 iovss.n1929 9.0005
R2991 iovss.n2160 iovss.n1929 9.0005
R2992 iovss.n2162 iovss.n1929 9.0005
R2993 iovss.n2241 iovss.n1929 9.0005
R2994 iovss.n1961 iovss.n1905 9.0005
R2995 iovss.n2095 iovss.n1905 9.0005
R2996 iovss.n2243 iovss.n1905 9.0005
R2997 iovss.n1905 iovss.n1891 9.0005
R2998 iovss.n1960 iovss.n1905 9.0005
R2999 iovss.n2098 iovss.n1905 9.0005
R3000 iovss.n1958 iovss.n1905 9.0005
R3001 iovss.n2101 iovss.n1905 9.0005
R3002 iovss.n1957 iovss.n1905 9.0005
R3003 iovss.n2104 iovss.n1905 9.0005
R3004 iovss.n1956 iovss.n1905 9.0005
R3005 iovss.n2106 iovss.n1905 9.0005
R3006 iovss.n1955 iovss.n1905 9.0005
R3007 iovss.n2109 iovss.n1905 9.0005
R3008 iovss.n1954 iovss.n1905 9.0005
R3009 iovss.n2111 iovss.n1905 9.0005
R3010 iovss.n1953 iovss.n1905 9.0005
R3011 iovss.n2114 iovss.n1905 9.0005
R3012 iovss.n1952 iovss.n1905 9.0005
R3013 iovss.n2116 iovss.n1905 9.0005
R3014 iovss.n1951 iovss.n1905 9.0005
R3015 iovss.n2119 iovss.n1905 9.0005
R3016 iovss.n1950 iovss.n1905 9.0005
R3017 iovss.n2121 iovss.n1905 9.0005
R3018 iovss.n1949 iovss.n1905 9.0005
R3019 iovss.n2124 iovss.n1905 9.0005
R3020 iovss.n1948 iovss.n1905 9.0005
R3021 iovss.n2126 iovss.n1905 9.0005
R3022 iovss.n1947 iovss.n1905 9.0005
R3023 iovss.n2129 iovss.n1905 9.0005
R3024 iovss.n1946 iovss.n1905 9.0005
R3025 iovss.n2131 iovss.n1905 9.0005
R3026 iovss.n1945 iovss.n1905 9.0005
R3027 iovss.n2160 iovss.n1905 9.0005
R3028 iovss.n2162 iovss.n1905 9.0005
R3029 iovss.n2241 iovss.n1905 9.0005
R3030 iovss.n1961 iovss.n1930 9.0005
R3031 iovss.n2095 iovss.n1930 9.0005
R3032 iovss.n2243 iovss.n1930 9.0005
R3033 iovss.n1930 iovss.n1891 9.0005
R3034 iovss.n1960 iovss.n1930 9.0005
R3035 iovss.n2098 iovss.n1930 9.0005
R3036 iovss.n1958 iovss.n1930 9.0005
R3037 iovss.n2101 iovss.n1930 9.0005
R3038 iovss.n1957 iovss.n1930 9.0005
R3039 iovss.n2104 iovss.n1930 9.0005
R3040 iovss.n1956 iovss.n1930 9.0005
R3041 iovss.n2106 iovss.n1930 9.0005
R3042 iovss.n1955 iovss.n1930 9.0005
R3043 iovss.n2109 iovss.n1930 9.0005
R3044 iovss.n1954 iovss.n1930 9.0005
R3045 iovss.n2111 iovss.n1930 9.0005
R3046 iovss.n1953 iovss.n1930 9.0005
R3047 iovss.n2114 iovss.n1930 9.0005
R3048 iovss.n1952 iovss.n1930 9.0005
R3049 iovss.n2116 iovss.n1930 9.0005
R3050 iovss.n1951 iovss.n1930 9.0005
R3051 iovss.n2119 iovss.n1930 9.0005
R3052 iovss.n1950 iovss.n1930 9.0005
R3053 iovss.n2121 iovss.n1930 9.0005
R3054 iovss.n1949 iovss.n1930 9.0005
R3055 iovss.n2124 iovss.n1930 9.0005
R3056 iovss.n1948 iovss.n1930 9.0005
R3057 iovss.n2126 iovss.n1930 9.0005
R3058 iovss.n1947 iovss.n1930 9.0005
R3059 iovss.n2129 iovss.n1930 9.0005
R3060 iovss.n1946 iovss.n1930 9.0005
R3061 iovss.n2131 iovss.n1930 9.0005
R3062 iovss.n1945 iovss.n1930 9.0005
R3063 iovss.n2160 iovss.n1930 9.0005
R3064 iovss.n2162 iovss.n1930 9.0005
R3065 iovss.n2241 iovss.n1930 9.0005
R3066 iovss.n1961 iovss.n1904 9.0005
R3067 iovss.n2095 iovss.n1904 9.0005
R3068 iovss.n2243 iovss.n1904 9.0005
R3069 iovss.n1904 iovss.n1891 9.0005
R3070 iovss.n1960 iovss.n1904 9.0005
R3071 iovss.n2098 iovss.n1904 9.0005
R3072 iovss.n1958 iovss.n1904 9.0005
R3073 iovss.n2101 iovss.n1904 9.0005
R3074 iovss.n1957 iovss.n1904 9.0005
R3075 iovss.n2104 iovss.n1904 9.0005
R3076 iovss.n1956 iovss.n1904 9.0005
R3077 iovss.n2106 iovss.n1904 9.0005
R3078 iovss.n1955 iovss.n1904 9.0005
R3079 iovss.n2109 iovss.n1904 9.0005
R3080 iovss.n1954 iovss.n1904 9.0005
R3081 iovss.n2111 iovss.n1904 9.0005
R3082 iovss.n1953 iovss.n1904 9.0005
R3083 iovss.n2114 iovss.n1904 9.0005
R3084 iovss.n1952 iovss.n1904 9.0005
R3085 iovss.n2116 iovss.n1904 9.0005
R3086 iovss.n1951 iovss.n1904 9.0005
R3087 iovss.n2119 iovss.n1904 9.0005
R3088 iovss.n1950 iovss.n1904 9.0005
R3089 iovss.n2121 iovss.n1904 9.0005
R3090 iovss.n1949 iovss.n1904 9.0005
R3091 iovss.n2124 iovss.n1904 9.0005
R3092 iovss.n1948 iovss.n1904 9.0005
R3093 iovss.n2126 iovss.n1904 9.0005
R3094 iovss.n1947 iovss.n1904 9.0005
R3095 iovss.n2129 iovss.n1904 9.0005
R3096 iovss.n1946 iovss.n1904 9.0005
R3097 iovss.n2131 iovss.n1904 9.0005
R3098 iovss.n1945 iovss.n1904 9.0005
R3099 iovss.n2160 iovss.n1904 9.0005
R3100 iovss.n2162 iovss.n1904 9.0005
R3101 iovss.n2241 iovss.n1904 9.0005
R3102 iovss.n1961 iovss.n1931 9.0005
R3103 iovss.n2095 iovss.n1931 9.0005
R3104 iovss.n2243 iovss.n1931 9.0005
R3105 iovss.n1931 iovss.n1891 9.0005
R3106 iovss.n1960 iovss.n1931 9.0005
R3107 iovss.n2098 iovss.n1931 9.0005
R3108 iovss.n1958 iovss.n1931 9.0005
R3109 iovss.n2101 iovss.n1931 9.0005
R3110 iovss.n1957 iovss.n1931 9.0005
R3111 iovss.n2104 iovss.n1931 9.0005
R3112 iovss.n1956 iovss.n1931 9.0005
R3113 iovss.n2106 iovss.n1931 9.0005
R3114 iovss.n1955 iovss.n1931 9.0005
R3115 iovss.n2109 iovss.n1931 9.0005
R3116 iovss.n1954 iovss.n1931 9.0005
R3117 iovss.n2111 iovss.n1931 9.0005
R3118 iovss.n1953 iovss.n1931 9.0005
R3119 iovss.n2114 iovss.n1931 9.0005
R3120 iovss.n1952 iovss.n1931 9.0005
R3121 iovss.n2116 iovss.n1931 9.0005
R3122 iovss.n1951 iovss.n1931 9.0005
R3123 iovss.n2119 iovss.n1931 9.0005
R3124 iovss.n1950 iovss.n1931 9.0005
R3125 iovss.n2121 iovss.n1931 9.0005
R3126 iovss.n1949 iovss.n1931 9.0005
R3127 iovss.n2124 iovss.n1931 9.0005
R3128 iovss.n1948 iovss.n1931 9.0005
R3129 iovss.n2126 iovss.n1931 9.0005
R3130 iovss.n1947 iovss.n1931 9.0005
R3131 iovss.n2129 iovss.n1931 9.0005
R3132 iovss.n1946 iovss.n1931 9.0005
R3133 iovss.n2131 iovss.n1931 9.0005
R3134 iovss.n1945 iovss.n1931 9.0005
R3135 iovss.n2160 iovss.n1931 9.0005
R3136 iovss.n2162 iovss.n1931 9.0005
R3137 iovss.n2241 iovss.n1931 9.0005
R3138 iovss.n1961 iovss.n1903 9.0005
R3139 iovss.n2095 iovss.n1903 9.0005
R3140 iovss.n2243 iovss.n1903 9.0005
R3141 iovss.n1903 iovss.n1891 9.0005
R3142 iovss.n1960 iovss.n1903 9.0005
R3143 iovss.n2098 iovss.n1903 9.0005
R3144 iovss.n1958 iovss.n1903 9.0005
R3145 iovss.n2101 iovss.n1903 9.0005
R3146 iovss.n1957 iovss.n1903 9.0005
R3147 iovss.n2104 iovss.n1903 9.0005
R3148 iovss.n1956 iovss.n1903 9.0005
R3149 iovss.n2106 iovss.n1903 9.0005
R3150 iovss.n1955 iovss.n1903 9.0005
R3151 iovss.n2109 iovss.n1903 9.0005
R3152 iovss.n1954 iovss.n1903 9.0005
R3153 iovss.n2111 iovss.n1903 9.0005
R3154 iovss.n1953 iovss.n1903 9.0005
R3155 iovss.n2114 iovss.n1903 9.0005
R3156 iovss.n1952 iovss.n1903 9.0005
R3157 iovss.n2116 iovss.n1903 9.0005
R3158 iovss.n1951 iovss.n1903 9.0005
R3159 iovss.n2119 iovss.n1903 9.0005
R3160 iovss.n1950 iovss.n1903 9.0005
R3161 iovss.n2121 iovss.n1903 9.0005
R3162 iovss.n1949 iovss.n1903 9.0005
R3163 iovss.n2124 iovss.n1903 9.0005
R3164 iovss.n1948 iovss.n1903 9.0005
R3165 iovss.n2126 iovss.n1903 9.0005
R3166 iovss.n1947 iovss.n1903 9.0005
R3167 iovss.n2129 iovss.n1903 9.0005
R3168 iovss.n1946 iovss.n1903 9.0005
R3169 iovss.n2131 iovss.n1903 9.0005
R3170 iovss.n1945 iovss.n1903 9.0005
R3171 iovss.n2160 iovss.n1903 9.0005
R3172 iovss.n2162 iovss.n1903 9.0005
R3173 iovss.n2241 iovss.n1903 9.0005
R3174 iovss.n1961 iovss.n1932 9.0005
R3175 iovss.n2095 iovss.n1932 9.0005
R3176 iovss.n2243 iovss.n1932 9.0005
R3177 iovss.n1932 iovss.n1891 9.0005
R3178 iovss.n1960 iovss.n1932 9.0005
R3179 iovss.n2098 iovss.n1932 9.0005
R3180 iovss.n1958 iovss.n1932 9.0005
R3181 iovss.n2101 iovss.n1932 9.0005
R3182 iovss.n1957 iovss.n1932 9.0005
R3183 iovss.n2104 iovss.n1932 9.0005
R3184 iovss.n1956 iovss.n1932 9.0005
R3185 iovss.n2106 iovss.n1932 9.0005
R3186 iovss.n1955 iovss.n1932 9.0005
R3187 iovss.n2109 iovss.n1932 9.0005
R3188 iovss.n1954 iovss.n1932 9.0005
R3189 iovss.n2111 iovss.n1932 9.0005
R3190 iovss.n1953 iovss.n1932 9.0005
R3191 iovss.n2114 iovss.n1932 9.0005
R3192 iovss.n1952 iovss.n1932 9.0005
R3193 iovss.n2116 iovss.n1932 9.0005
R3194 iovss.n1951 iovss.n1932 9.0005
R3195 iovss.n2119 iovss.n1932 9.0005
R3196 iovss.n1950 iovss.n1932 9.0005
R3197 iovss.n2121 iovss.n1932 9.0005
R3198 iovss.n1949 iovss.n1932 9.0005
R3199 iovss.n2124 iovss.n1932 9.0005
R3200 iovss.n1948 iovss.n1932 9.0005
R3201 iovss.n2126 iovss.n1932 9.0005
R3202 iovss.n1947 iovss.n1932 9.0005
R3203 iovss.n2129 iovss.n1932 9.0005
R3204 iovss.n1946 iovss.n1932 9.0005
R3205 iovss.n2131 iovss.n1932 9.0005
R3206 iovss.n1945 iovss.n1932 9.0005
R3207 iovss.n2160 iovss.n1932 9.0005
R3208 iovss.n2162 iovss.n1932 9.0005
R3209 iovss.n2241 iovss.n1932 9.0005
R3210 iovss.n1961 iovss.n1902 9.0005
R3211 iovss.n2095 iovss.n1902 9.0005
R3212 iovss.n2243 iovss.n1902 9.0005
R3213 iovss.n1902 iovss.n1891 9.0005
R3214 iovss.n1960 iovss.n1902 9.0005
R3215 iovss.n2098 iovss.n1902 9.0005
R3216 iovss.n1958 iovss.n1902 9.0005
R3217 iovss.n2101 iovss.n1902 9.0005
R3218 iovss.n1957 iovss.n1902 9.0005
R3219 iovss.n2104 iovss.n1902 9.0005
R3220 iovss.n1956 iovss.n1902 9.0005
R3221 iovss.n2106 iovss.n1902 9.0005
R3222 iovss.n1955 iovss.n1902 9.0005
R3223 iovss.n2109 iovss.n1902 9.0005
R3224 iovss.n1954 iovss.n1902 9.0005
R3225 iovss.n2111 iovss.n1902 9.0005
R3226 iovss.n1953 iovss.n1902 9.0005
R3227 iovss.n2114 iovss.n1902 9.0005
R3228 iovss.n1952 iovss.n1902 9.0005
R3229 iovss.n2116 iovss.n1902 9.0005
R3230 iovss.n1951 iovss.n1902 9.0005
R3231 iovss.n2119 iovss.n1902 9.0005
R3232 iovss.n1950 iovss.n1902 9.0005
R3233 iovss.n2121 iovss.n1902 9.0005
R3234 iovss.n1949 iovss.n1902 9.0005
R3235 iovss.n2124 iovss.n1902 9.0005
R3236 iovss.n1948 iovss.n1902 9.0005
R3237 iovss.n2126 iovss.n1902 9.0005
R3238 iovss.n1947 iovss.n1902 9.0005
R3239 iovss.n2129 iovss.n1902 9.0005
R3240 iovss.n1946 iovss.n1902 9.0005
R3241 iovss.n2131 iovss.n1902 9.0005
R3242 iovss.n1945 iovss.n1902 9.0005
R3243 iovss.n2160 iovss.n1902 9.0005
R3244 iovss.n2162 iovss.n1902 9.0005
R3245 iovss.n2241 iovss.n1902 9.0005
R3246 iovss.n1961 iovss.n1933 9.0005
R3247 iovss.n2095 iovss.n1933 9.0005
R3248 iovss.n2243 iovss.n1933 9.0005
R3249 iovss.n1933 iovss.n1891 9.0005
R3250 iovss.n1960 iovss.n1933 9.0005
R3251 iovss.n2098 iovss.n1933 9.0005
R3252 iovss.n1958 iovss.n1933 9.0005
R3253 iovss.n2101 iovss.n1933 9.0005
R3254 iovss.n1957 iovss.n1933 9.0005
R3255 iovss.n2104 iovss.n1933 9.0005
R3256 iovss.n1956 iovss.n1933 9.0005
R3257 iovss.n2106 iovss.n1933 9.0005
R3258 iovss.n1955 iovss.n1933 9.0005
R3259 iovss.n2109 iovss.n1933 9.0005
R3260 iovss.n1954 iovss.n1933 9.0005
R3261 iovss.n2111 iovss.n1933 9.0005
R3262 iovss.n1953 iovss.n1933 9.0005
R3263 iovss.n2114 iovss.n1933 9.0005
R3264 iovss.n1952 iovss.n1933 9.0005
R3265 iovss.n2116 iovss.n1933 9.0005
R3266 iovss.n1951 iovss.n1933 9.0005
R3267 iovss.n2119 iovss.n1933 9.0005
R3268 iovss.n1950 iovss.n1933 9.0005
R3269 iovss.n2121 iovss.n1933 9.0005
R3270 iovss.n1949 iovss.n1933 9.0005
R3271 iovss.n2124 iovss.n1933 9.0005
R3272 iovss.n1948 iovss.n1933 9.0005
R3273 iovss.n2126 iovss.n1933 9.0005
R3274 iovss.n1947 iovss.n1933 9.0005
R3275 iovss.n2129 iovss.n1933 9.0005
R3276 iovss.n1946 iovss.n1933 9.0005
R3277 iovss.n2131 iovss.n1933 9.0005
R3278 iovss.n1945 iovss.n1933 9.0005
R3279 iovss.n2160 iovss.n1933 9.0005
R3280 iovss.n2162 iovss.n1933 9.0005
R3281 iovss.n2241 iovss.n1933 9.0005
R3282 iovss.n1961 iovss.n1901 9.0005
R3283 iovss.n2095 iovss.n1901 9.0005
R3284 iovss.n2243 iovss.n1901 9.0005
R3285 iovss.n1901 iovss.n1891 9.0005
R3286 iovss.n1960 iovss.n1901 9.0005
R3287 iovss.n2098 iovss.n1901 9.0005
R3288 iovss.n1958 iovss.n1901 9.0005
R3289 iovss.n2101 iovss.n1901 9.0005
R3290 iovss.n1957 iovss.n1901 9.0005
R3291 iovss.n2104 iovss.n1901 9.0005
R3292 iovss.n1956 iovss.n1901 9.0005
R3293 iovss.n2106 iovss.n1901 9.0005
R3294 iovss.n1955 iovss.n1901 9.0005
R3295 iovss.n2109 iovss.n1901 9.0005
R3296 iovss.n1954 iovss.n1901 9.0005
R3297 iovss.n2111 iovss.n1901 9.0005
R3298 iovss.n1953 iovss.n1901 9.0005
R3299 iovss.n2114 iovss.n1901 9.0005
R3300 iovss.n1952 iovss.n1901 9.0005
R3301 iovss.n2116 iovss.n1901 9.0005
R3302 iovss.n1951 iovss.n1901 9.0005
R3303 iovss.n2119 iovss.n1901 9.0005
R3304 iovss.n1950 iovss.n1901 9.0005
R3305 iovss.n2121 iovss.n1901 9.0005
R3306 iovss.n1949 iovss.n1901 9.0005
R3307 iovss.n2124 iovss.n1901 9.0005
R3308 iovss.n1948 iovss.n1901 9.0005
R3309 iovss.n2126 iovss.n1901 9.0005
R3310 iovss.n1947 iovss.n1901 9.0005
R3311 iovss.n2129 iovss.n1901 9.0005
R3312 iovss.n1946 iovss.n1901 9.0005
R3313 iovss.n2131 iovss.n1901 9.0005
R3314 iovss.n1945 iovss.n1901 9.0005
R3315 iovss.n2160 iovss.n1901 9.0005
R3316 iovss.n2162 iovss.n1901 9.0005
R3317 iovss.n2241 iovss.n1901 9.0005
R3318 iovss.n1961 iovss.n1934 9.0005
R3319 iovss.n2095 iovss.n1934 9.0005
R3320 iovss.n2243 iovss.n1934 9.0005
R3321 iovss.n1934 iovss.n1891 9.0005
R3322 iovss.n1960 iovss.n1934 9.0005
R3323 iovss.n2098 iovss.n1934 9.0005
R3324 iovss.n1958 iovss.n1934 9.0005
R3325 iovss.n2101 iovss.n1934 9.0005
R3326 iovss.n1957 iovss.n1934 9.0005
R3327 iovss.n2104 iovss.n1934 9.0005
R3328 iovss.n1956 iovss.n1934 9.0005
R3329 iovss.n2106 iovss.n1934 9.0005
R3330 iovss.n1955 iovss.n1934 9.0005
R3331 iovss.n2109 iovss.n1934 9.0005
R3332 iovss.n1954 iovss.n1934 9.0005
R3333 iovss.n2111 iovss.n1934 9.0005
R3334 iovss.n1953 iovss.n1934 9.0005
R3335 iovss.n2114 iovss.n1934 9.0005
R3336 iovss.n1952 iovss.n1934 9.0005
R3337 iovss.n2116 iovss.n1934 9.0005
R3338 iovss.n1951 iovss.n1934 9.0005
R3339 iovss.n2119 iovss.n1934 9.0005
R3340 iovss.n1950 iovss.n1934 9.0005
R3341 iovss.n2121 iovss.n1934 9.0005
R3342 iovss.n1949 iovss.n1934 9.0005
R3343 iovss.n2124 iovss.n1934 9.0005
R3344 iovss.n1948 iovss.n1934 9.0005
R3345 iovss.n2126 iovss.n1934 9.0005
R3346 iovss.n1947 iovss.n1934 9.0005
R3347 iovss.n2129 iovss.n1934 9.0005
R3348 iovss.n1946 iovss.n1934 9.0005
R3349 iovss.n2131 iovss.n1934 9.0005
R3350 iovss.n1945 iovss.n1934 9.0005
R3351 iovss.n2160 iovss.n1934 9.0005
R3352 iovss.n2162 iovss.n1934 9.0005
R3353 iovss.n2241 iovss.n1934 9.0005
R3354 iovss.n1961 iovss.n1900 9.0005
R3355 iovss.n2095 iovss.n1900 9.0005
R3356 iovss.n2243 iovss.n1900 9.0005
R3357 iovss.n1900 iovss.n1891 9.0005
R3358 iovss.n1960 iovss.n1900 9.0005
R3359 iovss.n2098 iovss.n1900 9.0005
R3360 iovss.n1958 iovss.n1900 9.0005
R3361 iovss.n2101 iovss.n1900 9.0005
R3362 iovss.n1957 iovss.n1900 9.0005
R3363 iovss.n2104 iovss.n1900 9.0005
R3364 iovss.n1956 iovss.n1900 9.0005
R3365 iovss.n2106 iovss.n1900 9.0005
R3366 iovss.n1955 iovss.n1900 9.0005
R3367 iovss.n2109 iovss.n1900 9.0005
R3368 iovss.n1954 iovss.n1900 9.0005
R3369 iovss.n2111 iovss.n1900 9.0005
R3370 iovss.n1953 iovss.n1900 9.0005
R3371 iovss.n2114 iovss.n1900 9.0005
R3372 iovss.n1952 iovss.n1900 9.0005
R3373 iovss.n2116 iovss.n1900 9.0005
R3374 iovss.n1951 iovss.n1900 9.0005
R3375 iovss.n2119 iovss.n1900 9.0005
R3376 iovss.n1950 iovss.n1900 9.0005
R3377 iovss.n2121 iovss.n1900 9.0005
R3378 iovss.n1949 iovss.n1900 9.0005
R3379 iovss.n2124 iovss.n1900 9.0005
R3380 iovss.n1948 iovss.n1900 9.0005
R3381 iovss.n2126 iovss.n1900 9.0005
R3382 iovss.n1947 iovss.n1900 9.0005
R3383 iovss.n2129 iovss.n1900 9.0005
R3384 iovss.n1946 iovss.n1900 9.0005
R3385 iovss.n2131 iovss.n1900 9.0005
R3386 iovss.n1945 iovss.n1900 9.0005
R3387 iovss.n2160 iovss.n1900 9.0005
R3388 iovss.n2162 iovss.n1900 9.0005
R3389 iovss.n2241 iovss.n1900 9.0005
R3390 iovss.n1961 iovss.n1935 9.0005
R3391 iovss.n2095 iovss.n1935 9.0005
R3392 iovss.n2243 iovss.n1935 9.0005
R3393 iovss.n1935 iovss.n1891 9.0005
R3394 iovss.n1960 iovss.n1935 9.0005
R3395 iovss.n2098 iovss.n1935 9.0005
R3396 iovss.n1958 iovss.n1935 9.0005
R3397 iovss.n2101 iovss.n1935 9.0005
R3398 iovss.n1957 iovss.n1935 9.0005
R3399 iovss.n2104 iovss.n1935 9.0005
R3400 iovss.n1956 iovss.n1935 9.0005
R3401 iovss.n2106 iovss.n1935 9.0005
R3402 iovss.n1955 iovss.n1935 9.0005
R3403 iovss.n2109 iovss.n1935 9.0005
R3404 iovss.n1954 iovss.n1935 9.0005
R3405 iovss.n2111 iovss.n1935 9.0005
R3406 iovss.n1953 iovss.n1935 9.0005
R3407 iovss.n2114 iovss.n1935 9.0005
R3408 iovss.n1952 iovss.n1935 9.0005
R3409 iovss.n2116 iovss.n1935 9.0005
R3410 iovss.n1951 iovss.n1935 9.0005
R3411 iovss.n2119 iovss.n1935 9.0005
R3412 iovss.n1950 iovss.n1935 9.0005
R3413 iovss.n2121 iovss.n1935 9.0005
R3414 iovss.n1949 iovss.n1935 9.0005
R3415 iovss.n2124 iovss.n1935 9.0005
R3416 iovss.n1948 iovss.n1935 9.0005
R3417 iovss.n2126 iovss.n1935 9.0005
R3418 iovss.n1947 iovss.n1935 9.0005
R3419 iovss.n2129 iovss.n1935 9.0005
R3420 iovss.n1946 iovss.n1935 9.0005
R3421 iovss.n2131 iovss.n1935 9.0005
R3422 iovss.n1945 iovss.n1935 9.0005
R3423 iovss.n2160 iovss.n1935 9.0005
R3424 iovss.n2162 iovss.n1935 9.0005
R3425 iovss.n2241 iovss.n1935 9.0005
R3426 iovss.n1961 iovss.n1899 9.0005
R3427 iovss.n2095 iovss.n1899 9.0005
R3428 iovss.n2243 iovss.n1899 9.0005
R3429 iovss.n1899 iovss.n1891 9.0005
R3430 iovss.n1960 iovss.n1899 9.0005
R3431 iovss.n2098 iovss.n1899 9.0005
R3432 iovss.n1958 iovss.n1899 9.0005
R3433 iovss.n2101 iovss.n1899 9.0005
R3434 iovss.n1957 iovss.n1899 9.0005
R3435 iovss.n2104 iovss.n1899 9.0005
R3436 iovss.n1956 iovss.n1899 9.0005
R3437 iovss.n2106 iovss.n1899 9.0005
R3438 iovss.n1955 iovss.n1899 9.0005
R3439 iovss.n2109 iovss.n1899 9.0005
R3440 iovss.n1954 iovss.n1899 9.0005
R3441 iovss.n2111 iovss.n1899 9.0005
R3442 iovss.n1953 iovss.n1899 9.0005
R3443 iovss.n2114 iovss.n1899 9.0005
R3444 iovss.n1952 iovss.n1899 9.0005
R3445 iovss.n2116 iovss.n1899 9.0005
R3446 iovss.n1951 iovss.n1899 9.0005
R3447 iovss.n2119 iovss.n1899 9.0005
R3448 iovss.n1950 iovss.n1899 9.0005
R3449 iovss.n2121 iovss.n1899 9.0005
R3450 iovss.n1949 iovss.n1899 9.0005
R3451 iovss.n2124 iovss.n1899 9.0005
R3452 iovss.n1948 iovss.n1899 9.0005
R3453 iovss.n2126 iovss.n1899 9.0005
R3454 iovss.n1947 iovss.n1899 9.0005
R3455 iovss.n2129 iovss.n1899 9.0005
R3456 iovss.n1946 iovss.n1899 9.0005
R3457 iovss.n2131 iovss.n1899 9.0005
R3458 iovss.n1945 iovss.n1899 9.0005
R3459 iovss.n2160 iovss.n1899 9.0005
R3460 iovss.n2162 iovss.n1899 9.0005
R3461 iovss.n2241 iovss.n1899 9.0005
R3462 iovss.n1961 iovss.n1936 9.0005
R3463 iovss.n2095 iovss.n1936 9.0005
R3464 iovss.n2243 iovss.n1936 9.0005
R3465 iovss.n1936 iovss.n1891 9.0005
R3466 iovss.n1960 iovss.n1936 9.0005
R3467 iovss.n2098 iovss.n1936 9.0005
R3468 iovss.n1958 iovss.n1936 9.0005
R3469 iovss.n2101 iovss.n1936 9.0005
R3470 iovss.n1957 iovss.n1936 9.0005
R3471 iovss.n2104 iovss.n1936 9.0005
R3472 iovss.n1956 iovss.n1936 9.0005
R3473 iovss.n2106 iovss.n1936 9.0005
R3474 iovss.n1955 iovss.n1936 9.0005
R3475 iovss.n2109 iovss.n1936 9.0005
R3476 iovss.n1954 iovss.n1936 9.0005
R3477 iovss.n2111 iovss.n1936 9.0005
R3478 iovss.n1953 iovss.n1936 9.0005
R3479 iovss.n2114 iovss.n1936 9.0005
R3480 iovss.n1952 iovss.n1936 9.0005
R3481 iovss.n2116 iovss.n1936 9.0005
R3482 iovss.n1951 iovss.n1936 9.0005
R3483 iovss.n2119 iovss.n1936 9.0005
R3484 iovss.n1950 iovss.n1936 9.0005
R3485 iovss.n2121 iovss.n1936 9.0005
R3486 iovss.n1949 iovss.n1936 9.0005
R3487 iovss.n2124 iovss.n1936 9.0005
R3488 iovss.n1948 iovss.n1936 9.0005
R3489 iovss.n2126 iovss.n1936 9.0005
R3490 iovss.n1947 iovss.n1936 9.0005
R3491 iovss.n2129 iovss.n1936 9.0005
R3492 iovss.n1946 iovss.n1936 9.0005
R3493 iovss.n2131 iovss.n1936 9.0005
R3494 iovss.n1945 iovss.n1936 9.0005
R3495 iovss.n2160 iovss.n1936 9.0005
R3496 iovss.n2162 iovss.n1936 9.0005
R3497 iovss.n2241 iovss.n1936 9.0005
R3498 iovss.n1961 iovss.n1898 9.0005
R3499 iovss.n2095 iovss.n1898 9.0005
R3500 iovss.n2243 iovss.n1898 9.0005
R3501 iovss.n1898 iovss.n1891 9.0005
R3502 iovss.n1960 iovss.n1898 9.0005
R3503 iovss.n2098 iovss.n1898 9.0005
R3504 iovss.n1958 iovss.n1898 9.0005
R3505 iovss.n2101 iovss.n1898 9.0005
R3506 iovss.n1957 iovss.n1898 9.0005
R3507 iovss.n2104 iovss.n1898 9.0005
R3508 iovss.n1956 iovss.n1898 9.0005
R3509 iovss.n2106 iovss.n1898 9.0005
R3510 iovss.n1955 iovss.n1898 9.0005
R3511 iovss.n2109 iovss.n1898 9.0005
R3512 iovss.n1954 iovss.n1898 9.0005
R3513 iovss.n2111 iovss.n1898 9.0005
R3514 iovss.n1953 iovss.n1898 9.0005
R3515 iovss.n2114 iovss.n1898 9.0005
R3516 iovss.n1952 iovss.n1898 9.0005
R3517 iovss.n2116 iovss.n1898 9.0005
R3518 iovss.n1951 iovss.n1898 9.0005
R3519 iovss.n2119 iovss.n1898 9.0005
R3520 iovss.n1950 iovss.n1898 9.0005
R3521 iovss.n2121 iovss.n1898 9.0005
R3522 iovss.n1949 iovss.n1898 9.0005
R3523 iovss.n2124 iovss.n1898 9.0005
R3524 iovss.n1948 iovss.n1898 9.0005
R3525 iovss.n2126 iovss.n1898 9.0005
R3526 iovss.n1947 iovss.n1898 9.0005
R3527 iovss.n2129 iovss.n1898 9.0005
R3528 iovss.n1946 iovss.n1898 9.0005
R3529 iovss.n2131 iovss.n1898 9.0005
R3530 iovss.n1945 iovss.n1898 9.0005
R3531 iovss.n2160 iovss.n1898 9.0005
R3532 iovss.n2162 iovss.n1898 9.0005
R3533 iovss.n2241 iovss.n1898 9.0005
R3534 iovss.n1961 iovss.n1937 9.0005
R3535 iovss.n2095 iovss.n1937 9.0005
R3536 iovss.n2243 iovss.n1937 9.0005
R3537 iovss.n1937 iovss.n1891 9.0005
R3538 iovss.n1960 iovss.n1937 9.0005
R3539 iovss.n2098 iovss.n1937 9.0005
R3540 iovss.n1958 iovss.n1937 9.0005
R3541 iovss.n2101 iovss.n1937 9.0005
R3542 iovss.n1957 iovss.n1937 9.0005
R3543 iovss.n2104 iovss.n1937 9.0005
R3544 iovss.n1956 iovss.n1937 9.0005
R3545 iovss.n2106 iovss.n1937 9.0005
R3546 iovss.n1955 iovss.n1937 9.0005
R3547 iovss.n2109 iovss.n1937 9.0005
R3548 iovss.n1954 iovss.n1937 9.0005
R3549 iovss.n2111 iovss.n1937 9.0005
R3550 iovss.n1953 iovss.n1937 9.0005
R3551 iovss.n2114 iovss.n1937 9.0005
R3552 iovss.n1952 iovss.n1937 9.0005
R3553 iovss.n2116 iovss.n1937 9.0005
R3554 iovss.n1951 iovss.n1937 9.0005
R3555 iovss.n2119 iovss.n1937 9.0005
R3556 iovss.n1950 iovss.n1937 9.0005
R3557 iovss.n2121 iovss.n1937 9.0005
R3558 iovss.n1949 iovss.n1937 9.0005
R3559 iovss.n2124 iovss.n1937 9.0005
R3560 iovss.n1948 iovss.n1937 9.0005
R3561 iovss.n2126 iovss.n1937 9.0005
R3562 iovss.n1947 iovss.n1937 9.0005
R3563 iovss.n2129 iovss.n1937 9.0005
R3564 iovss.n1946 iovss.n1937 9.0005
R3565 iovss.n2131 iovss.n1937 9.0005
R3566 iovss.n1945 iovss.n1937 9.0005
R3567 iovss.n2160 iovss.n1937 9.0005
R3568 iovss.n2162 iovss.n1937 9.0005
R3569 iovss.n2241 iovss.n1937 9.0005
R3570 iovss.n1961 iovss.n1897 9.0005
R3571 iovss.n2095 iovss.n1897 9.0005
R3572 iovss.n2243 iovss.n1897 9.0005
R3573 iovss.n1897 iovss.n1891 9.0005
R3574 iovss.n1960 iovss.n1897 9.0005
R3575 iovss.n2098 iovss.n1897 9.0005
R3576 iovss.n1958 iovss.n1897 9.0005
R3577 iovss.n2101 iovss.n1897 9.0005
R3578 iovss.n1957 iovss.n1897 9.0005
R3579 iovss.n2104 iovss.n1897 9.0005
R3580 iovss.n1956 iovss.n1897 9.0005
R3581 iovss.n2106 iovss.n1897 9.0005
R3582 iovss.n1955 iovss.n1897 9.0005
R3583 iovss.n2109 iovss.n1897 9.0005
R3584 iovss.n1954 iovss.n1897 9.0005
R3585 iovss.n2111 iovss.n1897 9.0005
R3586 iovss.n1953 iovss.n1897 9.0005
R3587 iovss.n2114 iovss.n1897 9.0005
R3588 iovss.n1952 iovss.n1897 9.0005
R3589 iovss.n2116 iovss.n1897 9.0005
R3590 iovss.n1951 iovss.n1897 9.0005
R3591 iovss.n2119 iovss.n1897 9.0005
R3592 iovss.n1950 iovss.n1897 9.0005
R3593 iovss.n2121 iovss.n1897 9.0005
R3594 iovss.n1949 iovss.n1897 9.0005
R3595 iovss.n2124 iovss.n1897 9.0005
R3596 iovss.n1948 iovss.n1897 9.0005
R3597 iovss.n2126 iovss.n1897 9.0005
R3598 iovss.n1947 iovss.n1897 9.0005
R3599 iovss.n2129 iovss.n1897 9.0005
R3600 iovss.n1946 iovss.n1897 9.0005
R3601 iovss.n2131 iovss.n1897 9.0005
R3602 iovss.n1945 iovss.n1897 9.0005
R3603 iovss.n2160 iovss.n1897 9.0005
R3604 iovss.n2162 iovss.n1897 9.0005
R3605 iovss.n2241 iovss.n1897 9.0005
R3606 iovss.n1961 iovss.n1938 9.0005
R3607 iovss.n2095 iovss.n1938 9.0005
R3608 iovss.n2243 iovss.n1938 9.0005
R3609 iovss.n1938 iovss.n1891 9.0005
R3610 iovss.n1960 iovss.n1938 9.0005
R3611 iovss.n2098 iovss.n1938 9.0005
R3612 iovss.n1958 iovss.n1938 9.0005
R3613 iovss.n2101 iovss.n1938 9.0005
R3614 iovss.n1957 iovss.n1938 9.0005
R3615 iovss.n2104 iovss.n1938 9.0005
R3616 iovss.n1956 iovss.n1938 9.0005
R3617 iovss.n2106 iovss.n1938 9.0005
R3618 iovss.n1955 iovss.n1938 9.0005
R3619 iovss.n2109 iovss.n1938 9.0005
R3620 iovss.n1954 iovss.n1938 9.0005
R3621 iovss.n2111 iovss.n1938 9.0005
R3622 iovss.n1953 iovss.n1938 9.0005
R3623 iovss.n2114 iovss.n1938 9.0005
R3624 iovss.n1952 iovss.n1938 9.0005
R3625 iovss.n2116 iovss.n1938 9.0005
R3626 iovss.n1951 iovss.n1938 9.0005
R3627 iovss.n2119 iovss.n1938 9.0005
R3628 iovss.n1950 iovss.n1938 9.0005
R3629 iovss.n2121 iovss.n1938 9.0005
R3630 iovss.n1949 iovss.n1938 9.0005
R3631 iovss.n2124 iovss.n1938 9.0005
R3632 iovss.n1948 iovss.n1938 9.0005
R3633 iovss.n2126 iovss.n1938 9.0005
R3634 iovss.n1947 iovss.n1938 9.0005
R3635 iovss.n2129 iovss.n1938 9.0005
R3636 iovss.n1946 iovss.n1938 9.0005
R3637 iovss.n2131 iovss.n1938 9.0005
R3638 iovss.n1945 iovss.n1938 9.0005
R3639 iovss.n2160 iovss.n1938 9.0005
R3640 iovss.n2162 iovss.n1938 9.0005
R3641 iovss.n2241 iovss.n1938 9.0005
R3642 iovss.n1961 iovss.n1896 9.0005
R3643 iovss.n2095 iovss.n1896 9.0005
R3644 iovss.n2243 iovss.n1896 9.0005
R3645 iovss.n1896 iovss.n1891 9.0005
R3646 iovss.n1960 iovss.n1896 9.0005
R3647 iovss.n2098 iovss.n1896 9.0005
R3648 iovss.n1958 iovss.n1896 9.0005
R3649 iovss.n2101 iovss.n1896 9.0005
R3650 iovss.n1957 iovss.n1896 9.0005
R3651 iovss.n2104 iovss.n1896 9.0005
R3652 iovss.n1956 iovss.n1896 9.0005
R3653 iovss.n2106 iovss.n1896 9.0005
R3654 iovss.n1955 iovss.n1896 9.0005
R3655 iovss.n2109 iovss.n1896 9.0005
R3656 iovss.n1954 iovss.n1896 9.0005
R3657 iovss.n2111 iovss.n1896 9.0005
R3658 iovss.n1953 iovss.n1896 9.0005
R3659 iovss.n2114 iovss.n1896 9.0005
R3660 iovss.n1952 iovss.n1896 9.0005
R3661 iovss.n2116 iovss.n1896 9.0005
R3662 iovss.n1951 iovss.n1896 9.0005
R3663 iovss.n2119 iovss.n1896 9.0005
R3664 iovss.n1950 iovss.n1896 9.0005
R3665 iovss.n2121 iovss.n1896 9.0005
R3666 iovss.n1949 iovss.n1896 9.0005
R3667 iovss.n2124 iovss.n1896 9.0005
R3668 iovss.n1948 iovss.n1896 9.0005
R3669 iovss.n2126 iovss.n1896 9.0005
R3670 iovss.n1947 iovss.n1896 9.0005
R3671 iovss.n2129 iovss.n1896 9.0005
R3672 iovss.n1946 iovss.n1896 9.0005
R3673 iovss.n2131 iovss.n1896 9.0005
R3674 iovss.n1945 iovss.n1896 9.0005
R3675 iovss.n2160 iovss.n1896 9.0005
R3676 iovss.n2162 iovss.n1896 9.0005
R3677 iovss.n2241 iovss.n1896 9.0005
R3678 iovss.n1961 iovss.n1939 9.0005
R3679 iovss.n2095 iovss.n1939 9.0005
R3680 iovss.n2243 iovss.n1939 9.0005
R3681 iovss.n1939 iovss.n1891 9.0005
R3682 iovss.n1960 iovss.n1939 9.0005
R3683 iovss.n2098 iovss.n1939 9.0005
R3684 iovss.n1958 iovss.n1939 9.0005
R3685 iovss.n2101 iovss.n1939 9.0005
R3686 iovss.n1957 iovss.n1939 9.0005
R3687 iovss.n2104 iovss.n1939 9.0005
R3688 iovss.n1956 iovss.n1939 9.0005
R3689 iovss.n2106 iovss.n1939 9.0005
R3690 iovss.n1955 iovss.n1939 9.0005
R3691 iovss.n2109 iovss.n1939 9.0005
R3692 iovss.n1954 iovss.n1939 9.0005
R3693 iovss.n2111 iovss.n1939 9.0005
R3694 iovss.n1953 iovss.n1939 9.0005
R3695 iovss.n2114 iovss.n1939 9.0005
R3696 iovss.n1952 iovss.n1939 9.0005
R3697 iovss.n2116 iovss.n1939 9.0005
R3698 iovss.n1951 iovss.n1939 9.0005
R3699 iovss.n2119 iovss.n1939 9.0005
R3700 iovss.n1950 iovss.n1939 9.0005
R3701 iovss.n2121 iovss.n1939 9.0005
R3702 iovss.n1949 iovss.n1939 9.0005
R3703 iovss.n2124 iovss.n1939 9.0005
R3704 iovss.n1948 iovss.n1939 9.0005
R3705 iovss.n2126 iovss.n1939 9.0005
R3706 iovss.n1947 iovss.n1939 9.0005
R3707 iovss.n2129 iovss.n1939 9.0005
R3708 iovss.n1946 iovss.n1939 9.0005
R3709 iovss.n2131 iovss.n1939 9.0005
R3710 iovss.n1945 iovss.n1939 9.0005
R3711 iovss.n2160 iovss.n1939 9.0005
R3712 iovss.n2162 iovss.n1939 9.0005
R3713 iovss.n2241 iovss.n1939 9.0005
R3714 iovss.n1961 iovss.n1895 9.0005
R3715 iovss.n2095 iovss.n1895 9.0005
R3716 iovss.n2243 iovss.n1895 9.0005
R3717 iovss.n1895 iovss.n1891 9.0005
R3718 iovss.n1960 iovss.n1895 9.0005
R3719 iovss.n2098 iovss.n1895 9.0005
R3720 iovss.n1958 iovss.n1895 9.0005
R3721 iovss.n2101 iovss.n1895 9.0005
R3722 iovss.n1957 iovss.n1895 9.0005
R3723 iovss.n2104 iovss.n1895 9.0005
R3724 iovss.n1956 iovss.n1895 9.0005
R3725 iovss.n2106 iovss.n1895 9.0005
R3726 iovss.n1955 iovss.n1895 9.0005
R3727 iovss.n2109 iovss.n1895 9.0005
R3728 iovss.n1954 iovss.n1895 9.0005
R3729 iovss.n2111 iovss.n1895 9.0005
R3730 iovss.n1953 iovss.n1895 9.0005
R3731 iovss.n2114 iovss.n1895 9.0005
R3732 iovss.n1952 iovss.n1895 9.0005
R3733 iovss.n2116 iovss.n1895 9.0005
R3734 iovss.n1951 iovss.n1895 9.0005
R3735 iovss.n2119 iovss.n1895 9.0005
R3736 iovss.n1950 iovss.n1895 9.0005
R3737 iovss.n2121 iovss.n1895 9.0005
R3738 iovss.n1949 iovss.n1895 9.0005
R3739 iovss.n2124 iovss.n1895 9.0005
R3740 iovss.n1948 iovss.n1895 9.0005
R3741 iovss.n2126 iovss.n1895 9.0005
R3742 iovss.n1947 iovss.n1895 9.0005
R3743 iovss.n2129 iovss.n1895 9.0005
R3744 iovss.n1946 iovss.n1895 9.0005
R3745 iovss.n2131 iovss.n1895 9.0005
R3746 iovss.n1945 iovss.n1895 9.0005
R3747 iovss.n2160 iovss.n1895 9.0005
R3748 iovss.n2162 iovss.n1895 9.0005
R3749 iovss.n2241 iovss.n1895 9.0005
R3750 iovss.n1961 iovss.n1940 9.0005
R3751 iovss.n2095 iovss.n1940 9.0005
R3752 iovss.n2243 iovss.n1940 9.0005
R3753 iovss.n1940 iovss.n1891 9.0005
R3754 iovss.n1960 iovss.n1940 9.0005
R3755 iovss.n2098 iovss.n1940 9.0005
R3756 iovss.n1958 iovss.n1940 9.0005
R3757 iovss.n2101 iovss.n1940 9.0005
R3758 iovss.n1957 iovss.n1940 9.0005
R3759 iovss.n2104 iovss.n1940 9.0005
R3760 iovss.n1956 iovss.n1940 9.0005
R3761 iovss.n2106 iovss.n1940 9.0005
R3762 iovss.n1955 iovss.n1940 9.0005
R3763 iovss.n2109 iovss.n1940 9.0005
R3764 iovss.n1954 iovss.n1940 9.0005
R3765 iovss.n2111 iovss.n1940 9.0005
R3766 iovss.n1953 iovss.n1940 9.0005
R3767 iovss.n2114 iovss.n1940 9.0005
R3768 iovss.n1952 iovss.n1940 9.0005
R3769 iovss.n2116 iovss.n1940 9.0005
R3770 iovss.n1951 iovss.n1940 9.0005
R3771 iovss.n2119 iovss.n1940 9.0005
R3772 iovss.n1950 iovss.n1940 9.0005
R3773 iovss.n2121 iovss.n1940 9.0005
R3774 iovss.n1949 iovss.n1940 9.0005
R3775 iovss.n2124 iovss.n1940 9.0005
R3776 iovss.n1948 iovss.n1940 9.0005
R3777 iovss.n2126 iovss.n1940 9.0005
R3778 iovss.n1947 iovss.n1940 9.0005
R3779 iovss.n2129 iovss.n1940 9.0005
R3780 iovss.n1946 iovss.n1940 9.0005
R3781 iovss.n2131 iovss.n1940 9.0005
R3782 iovss.n1945 iovss.n1940 9.0005
R3783 iovss.n2160 iovss.n1940 9.0005
R3784 iovss.n2162 iovss.n1940 9.0005
R3785 iovss.n2241 iovss.n1940 9.0005
R3786 iovss.n1961 iovss.n1894 9.0005
R3787 iovss.n2095 iovss.n1894 9.0005
R3788 iovss.n2243 iovss.n1894 9.0005
R3789 iovss.n1894 iovss.n1891 9.0005
R3790 iovss.n1960 iovss.n1894 9.0005
R3791 iovss.n2098 iovss.n1894 9.0005
R3792 iovss.n1958 iovss.n1894 9.0005
R3793 iovss.n2101 iovss.n1894 9.0005
R3794 iovss.n1957 iovss.n1894 9.0005
R3795 iovss.n2104 iovss.n1894 9.0005
R3796 iovss.n1956 iovss.n1894 9.0005
R3797 iovss.n2106 iovss.n1894 9.0005
R3798 iovss.n1955 iovss.n1894 9.0005
R3799 iovss.n2109 iovss.n1894 9.0005
R3800 iovss.n1954 iovss.n1894 9.0005
R3801 iovss.n2111 iovss.n1894 9.0005
R3802 iovss.n1953 iovss.n1894 9.0005
R3803 iovss.n2114 iovss.n1894 9.0005
R3804 iovss.n1952 iovss.n1894 9.0005
R3805 iovss.n2116 iovss.n1894 9.0005
R3806 iovss.n1951 iovss.n1894 9.0005
R3807 iovss.n2119 iovss.n1894 9.0005
R3808 iovss.n1950 iovss.n1894 9.0005
R3809 iovss.n2121 iovss.n1894 9.0005
R3810 iovss.n1949 iovss.n1894 9.0005
R3811 iovss.n2124 iovss.n1894 9.0005
R3812 iovss.n1948 iovss.n1894 9.0005
R3813 iovss.n2126 iovss.n1894 9.0005
R3814 iovss.n1947 iovss.n1894 9.0005
R3815 iovss.n2129 iovss.n1894 9.0005
R3816 iovss.n1946 iovss.n1894 9.0005
R3817 iovss.n2131 iovss.n1894 9.0005
R3818 iovss.n1945 iovss.n1894 9.0005
R3819 iovss.n2160 iovss.n1894 9.0005
R3820 iovss.n2162 iovss.n1894 9.0005
R3821 iovss.n2241 iovss.n1894 9.0005
R3822 iovss.n1961 iovss.n1941 9.0005
R3823 iovss.n2095 iovss.n1941 9.0005
R3824 iovss.n2243 iovss.n1941 9.0005
R3825 iovss.n1941 iovss.n1891 9.0005
R3826 iovss.n1960 iovss.n1941 9.0005
R3827 iovss.n2098 iovss.n1941 9.0005
R3828 iovss.n1958 iovss.n1941 9.0005
R3829 iovss.n2101 iovss.n1941 9.0005
R3830 iovss.n1957 iovss.n1941 9.0005
R3831 iovss.n2104 iovss.n1941 9.0005
R3832 iovss.n1956 iovss.n1941 9.0005
R3833 iovss.n2106 iovss.n1941 9.0005
R3834 iovss.n1955 iovss.n1941 9.0005
R3835 iovss.n2109 iovss.n1941 9.0005
R3836 iovss.n1954 iovss.n1941 9.0005
R3837 iovss.n2111 iovss.n1941 9.0005
R3838 iovss.n1953 iovss.n1941 9.0005
R3839 iovss.n2114 iovss.n1941 9.0005
R3840 iovss.n1952 iovss.n1941 9.0005
R3841 iovss.n2116 iovss.n1941 9.0005
R3842 iovss.n1951 iovss.n1941 9.0005
R3843 iovss.n2119 iovss.n1941 9.0005
R3844 iovss.n1950 iovss.n1941 9.0005
R3845 iovss.n2121 iovss.n1941 9.0005
R3846 iovss.n1949 iovss.n1941 9.0005
R3847 iovss.n2124 iovss.n1941 9.0005
R3848 iovss.n1948 iovss.n1941 9.0005
R3849 iovss.n2126 iovss.n1941 9.0005
R3850 iovss.n1947 iovss.n1941 9.0005
R3851 iovss.n2129 iovss.n1941 9.0005
R3852 iovss.n1946 iovss.n1941 9.0005
R3853 iovss.n2131 iovss.n1941 9.0005
R3854 iovss.n1945 iovss.n1941 9.0005
R3855 iovss.n2160 iovss.n1941 9.0005
R3856 iovss.n2162 iovss.n1941 9.0005
R3857 iovss.n2241 iovss.n1941 9.0005
R3858 iovss.n1961 iovss.n1893 9.0005
R3859 iovss.n2095 iovss.n1893 9.0005
R3860 iovss.n2243 iovss.n1893 9.0005
R3861 iovss.n1893 iovss.n1891 9.0005
R3862 iovss.n1960 iovss.n1893 9.0005
R3863 iovss.n2098 iovss.n1893 9.0005
R3864 iovss.n1958 iovss.n1893 9.0005
R3865 iovss.n2101 iovss.n1893 9.0005
R3866 iovss.n1957 iovss.n1893 9.0005
R3867 iovss.n2104 iovss.n1893 9.0005
R3868 iovss.n1956 iovss.n1893 9.0005
R3869 iovss.n2106 iovss.n1893 9.0005
R3870 iovss.n1955 iovss.n1893 9.0005
R3871 iovss.n2109 iovss.n1893 9.0005
R3872 iovss.n1954 iovss.n1893 9.0005
R3873 iovss.n2111 iovss.n1893 9.0005
R3874 iovss.n1953 iovss.n1893 9.0005
R3875 iovss.n2114 iovss.n1893 9.0005
R3876 iovss.n1952 iovss.n1893 9.0005
R3877 iovss.n2116 iovss.n1893 9.0005
R3878 iovss.n1951 iovss.n1893 9.0005
R3879 iovss.n2119 iovss.n1893 9.0005
R3880 iovss.n1950 iovss.n1893 9.0005
R3881 iovss.n2121 iovss.n1893 9.0005
R3882 iovss.n1949 iovss.n1893 9.0005
R3883 iovss.n2124 iovss.n1893 9.0005
R3884 iovss.n1948 iovss.n1893 9.0005
R3885 iovss.n2126 iovss.n1893 9.0005
R3886 iovss.n1947 iovss.n1893 9.0005
R3887 iovss.n2129 iovss.n1893 9.0005
R3888 iovss.n1946 iovss.n1893 9.0005
R3889 iovss.n2131 iovss.n1893 9.0005
R3890 iovss.n1945 iovss.n1893 9.0005
R3891 iovss.n2160 iovss.n1893 9.0005
R3892 iovss.n2162 iovss.n1893 9.0005
R3893 iovss.n2241 iovss.n1893 9.0005
R3894 iovss.n1961 iovss.n1942 9.0005
R3895 iovss.n2095 iovss.n1942 9.0005
R3896 iovss.n2243 iovss.n1942 9.0005
R3897 iovss.n1942 iovss.n1891 9.0005
R3898 iovss.n1960 iovss.n1942 9.0005
R3899 iovss.n2098 iovss.n1942 9.0005
R3900 iovss.n1958 iovss.n1942 9.0005
R3901 iovss.n2101 iovss.n1942 9.0005
R3902 iovss.n1957 iovss.n1942 9.0005
R3903 iovss.n2104 iovss.n1942 9.0005
R3904 iovss.n1956 iovss.n1942 9.0005
R3905 iovss.n2106 iovss.n1942 9.0005
R3906 iovss.n1955 iovss.n1942 9.0005
R3907 iovss.n2109 iovss.n1942 9.0005
R3908 iovss.n1954 iovss.n1942 9.0005
R3909 iovss.n2111 iovss.n1942 9.0005
R3910 iovss.n1953 iovss.n1942 9.0005
R3911 iovss.n2114 iovss.n1942 9.0005
R3912 iovss.n1952 iovss.n1942 9.0005
R3913 iovss.n2116 iovss.n1942 9.0005
R3914 iovss.n1951 iovss.n1942 9.0005
R3915 iovss.n2119 iovss.n1942 9.0005
R3916 iovss.n1950 iovss.n1942 9.0005
R3917 iovss.n2121 iovss.n1942 9.0005
R3918 iovss.n1949 iovss.n1942 9.0005
R3919 iovss.n2124 iovss.n1942 9.0005
R3920 iovss.n1948 iovss.n1942 9.0005
R3921 iovss.n2126 iovss.n1942 9.0005
R3922 iovss.n1947 iovss.n1942 9.0005
R3923 iovss.n2129 iovss.n1942 9.0005
R3924 iovss.n1946 iovss.n1942 9.0005
R3925 iovss.n2131 iovss.n1942 9.0005
R3926 iovss.n1945 iovss.n1942 9.0005
R3927 iovss.n2160 iovss.n1942 9.0005
R3928 iovss.n2162 iovss.n1942 9.0005
R3929 iovss.n2241 iovss.n1942 9.0005
R3930 iovss.n1961 iovss.n1892 9.0005
R3931 iovss.n2095 iovss.n1892 9.0005
R3932 iovss.n2243 iovss.n1892 9.0005
R3933 iovss.n1892 iovss.n1891 9.0005
R3934 iovss.n1960 iovss.n1892 9.0005
R3935 iovss.n2098 iovss.n1892 9.0005
R3936 iovss.n1958 iovss.n1892 9.0005
R3937 iovss.n2101 iovss.n1892 9.0005
R3938 iovss.n1957 iovss.n1892 9.0005
R3939 iovss.n2104 iovss.n1892 9.0005
R3940 iovss.n1956 iovss.n1892 9.0005
R3941 iovss.n2106 iovss.n1892 9.0005
R3942 iovss.n1955 iovss.n1892 9.0005
R3943 iovss.n2109 iovss.n1892 9.0005
R3944 iovss.n1954 iovss.n1892 9.0005
R3945 iovss.n2111 iovss.n1892 9.0005
R3946 iovss.n1953 iovss.n1892 9.0005
R3947 iovss.n2114 iovss.n1892 9.0005
R3948 iovss.n1952 iovss.n1892 9.0005
R3949 iovss.n2116 iovss.n1892 9.0005
R3950 iovss.n1951 iovss.n1892 9.0005
R3951 iovss.n2119 iovss.n1892 9.0005
R3952 iovss.n1950 iovss.n1892 9.0005
R3953 iovss.n2121 iovss.n1892 9.0005
R3954 iovss.n1949 iovss.n1892 9.0005
R3955 iovss.n2124 iovss.n1892 9.0005
R3956 iovss.n1948 iovss.n1892 9.0005
R3957 iovss.n2126 iovss.n1892 9.0005
R3958 iovss.n1947 iovss.n1892 9.0005
R3959 iovss.n2129 iovss.n1892 9.0005
R3960 iovss.n1946 iovss.n1892 9.0005
R3961 iovss.n2131 iovss.n1892 9.0005
R3962 iovss.n1945 iovss.n1892 9.0005
R3963 iovss.n2160 iovss.n1892 9.0005
R3964 iovss.n2162 iovss.n1892 9.0005
R3965 iovss.n2241 iovss.n1892 9.0005
R3966 iovss.n2242 iovss.n1961 9.0005
R3967 iovss.n2242 iovss.n2095 9.0005
R3968 iovss.n2243 iovss.n2242 9.0005
R3969 iovss.n2242 iovss.n1891 9.0005
R3970 iovss.n2242 iovss.n1960 9.0005
R3971 iovss.n2242 iovss.n2098 9.0005
R3972 iovss.n2242 iovss.n1958 9.0005
R3973 iovss.n2242 iovss.n2101 9.0005
R3974 iovss.n2242 iovss.n1957 9.0005
R3975 iovss.n2242 iovss.n2104 9.0005
R3976 iovss.n2242 iovss.n1956 9.0005
R3977 iovss.n2242 iovss.n2106 9.0005
R3978 iovss.n2242 iovss.n1955 9.0005
R3979 iovss.n2242 iovss.n2109 9.0005
R3980 iovss.n2242 iovss.n1954 9.0005
R3981 iovss.n2242 iovss.n2111 9.0005
R3982 iovss.n2242 iovss.n1953 9.0005
R3983 iovss.n2242 iovss.n2114 9.0005
R3984 iovss.n2242 iovss.n1952 9.0005
R3985 iovss.n2242 iovss.n2116 9.0005
R3986 iovss.n2242 iovss.n1951 9.0005
R3987 iovss.n2242 iovss.n2119 9.0005
R3988 iovss.n2242 iovss.n1950 9.0005
R3989 iovss.n2242 iovss.n2121 9.0005
R3990 iovss.n2242 iovss.n1949 9.0005
R3991 iovss.n2242 iovss.n2124 9.0005
R3992 iovss.n2242 iovss.n1948 9.0005
R3993 iovss.n2242 iovss.n2126 9.0005
R3994 iovss.n2242 iovss.n1947 9.0005
R3995 iovss.n2242 iovss.n2129 9.0005
R3996 iovss.n2242 iovss.n1946 9.0005
R3997 iovss.n2242 iovss.n2131 9.0005
R3998 iovss.n2242 iovss.n1945 9.0005
R3999 iovss.n2242 iovss.n2160 9.0005
R4000 iovss.n2242 iovss.n2241 9.0005
R4001 iovss.n3079 iovss.n2925 9.0005
R4002 iovss.n3079 iovss.n2926 9.0005
R4003 iovss.n3072 iovss.n2929 9.0005
R4004 iovss.n2936 iovss.n2929 9.0005
R4005 iovss.n2982 iovss.n2929 9.0005
R4006 iovss.n2984 iovss.n2929 9.0005
R4007 iovss.n2986 iovss.n2929 9.0005
R4008 iovss.n2988 iovss.n2929 9.0005
R4009 iovss.n2990 iovss.n2929 9.0005
R4010 iovss.n2992 iovss.n2929 9.0005
R4011 iovss.n2994 iovss.n2929 9.0005
R4012 iovss.n2996 iovss.n2929 9.0005
R4013 iovss.n2998 iovss.n2929 9.0005
R4014 iovss.n3000 iovss.n2929 9.0005
R4015 iovss.n3002 iovss.n2929 9.0005
R4016 iovss.n3004 iovss.n2929 9.0005
R4017 iovss.n3006 iovss.n2929 9.0005
R4018 iovss.n3008 iovss.n2929 9.0005
R4019 iovss.n3010 iovss.n2929 9.0005
R4020 iovss.n3012 iovss.n2929 9.0005
R4021 iovss.n3014 iovss.n2929 9.0005
R4022 iovss.n3016 iovss.n2929 9.0005
R4023 iovss.n3018 iovss.n2929 9.0005
R4024 iovss.n3020 iovss.n2929 9.0005
R4025 iovss.n3022 iovss.n2929 9.0005
R4026 iovss.n3024 iovss.n2929 9.0005
R4027 iovss.n3026 iovss.n2929 9.0005
R4028 iovss.n3028 iovss.n2929 9.0005
R4029 iovss.n3030 iovss.n2929 9.0005
R4030 iovss.n3032 iovss.n2929 9.0005
R4031 iovss.n3034 iovss.n2929 9.0005
R4032 iovss.n3036 iovss.n2929 9.0005
R4033 iovss.n3038 iovss.n2929 9.0005
R4034 iovss.n3040 iovss.n2929 9.0005
R4035 iovss.n3042 iovss.n2929 9.0005
R4036 iovss.n3044 iovss.n2929 9.0005
R4037 iovss.n3046 iovss.n2929 9.0005
R4038 iovss.n3048 iovss.n2929 9.0005
R4039 iovss.n3050 iovss.n2929 9.0005
R4040 iovss.n3052 iovss.n2929 9.0005
R4041 iovss.n3054 iovss.n2929 9.0005
R4042 iovss.n3056 iovss.n2929 9.0005
R4043 iovss.n3058 iovss.n2929 9.0005
R4044 iovss.n3060 iovss.n2929 9.0005
R4045 iovss.n3062 iovss.n2929 9.0005
R4046 iovss.n3064 iovss.n2929 9.0005
R4047 iovss.n3066 iovss.n2929 9.0005
R4048 iovss.n3070 iovss.n3069 9.0005
R4049 iovss.n3069 iovss.n2929 9.0005
R4050 iovss.n3078 iovss.n2929 9.0005
R4051 iovss.n3076 iovss.n2929 9.0005
R4052 iovss.n3079 iovss.n3078 9.0005
R4053 iovss.n3098 iovss.n1138 9.0005
R4054 iovss.n3098 iovss.n1141 9.0005
R4055 iovss.n3095 iovss.n1141 9.0005
R4056 iovss.n3098 iovss.n1136 9.0005
R4057 iovss.n3095 iovss.n1136 9.0005
R4058 iovss.n3095 iovss.n3085 9.0005
R4059 iovss.n1218 iovss.n1115 9.0005
R4060 iovss.n3095 iovss.n1218 9.0005
R4061 iovss.n3098 iovss.n1144 9.0005
R4062 iovss.n3095 iovss.n1144 9.0005
R4063 iovss.n3098 iovss.n1135 9.0005
R4064 iovss.n3095 iovss.n1135 9.0005
R4065 iovss.n3098 iovss.n1147 9.0005
R4066 iovss.n3095 iovss.n1147 9.0005
R4067 iovss.n3098 iovss.n1134 9.0005
R4068 iovss.n3095 iovss.n1134 9.0005
R4069 iovss.n3098 iovss.n1150 9.0005
R4070 iovss.n3095 iovss.n1150 9.0005
R4071 iovss.n3098 iovss.n1133 9.0005
R4072 iovss.n3095 iovss.n1133 9.0005
R4073 iovss.n3098 iovss.n1153 9.0005
R4074 iovss.n3095 iovss.n1153 9.0005
R4075 iovss.n3098 iovss.n1132 9.0005
R4076 iovss.n3095 iovss.n1132 9.0005
R4077 iovss.n3098 iovss.n1155 9.0005
R4078 iovss.n3095 iovss.n1155 9.0005
R4079 iovss.n3095 iovss.n1216 9.0005
R4080 iovss.n3087 iovss.n1115 9.0005
R4081 iovss.n3095 iovss.n3087 9.0005
R4082 iovss.n3098 iovss.n1130 9.0005
R4083 iovss.n3095 iovss.n1130 9.0005
R4084 iovss.n3098 iovss.n1158 9.0005
R4085 iovss.n3095 iovss.n1158 9.0005
R4086 iovss.n3098 iovss.n1129 9.0005
R4087 iovss.n3095 iovss.n1129 9.0005
R4088 iovss.n3098 iovss.n1161 9.0005
R4089 iovss.n3095 iovss.n1161 9.0005
R4090 iovss.n3098 iovss.n1128 9.0005
R4091 iovss.n3095 iovss.n1128 9.0005
R4092 iovss.n3095 iovss.n3089 9.0005
R4093 iovss.n1214 iovss.n1115 9.0005
R4094 iovss.n3095 iovss.n1214 9.0005
R4095 iovss.n3098 iovss.n1164 9.0005
R4096 iovss.n3095 iovss.n1164 9.0005
R4097 iovss.n3098 iovss.n1127 9.0005
R4098 iovss.n3095 iovss.n1127 9.0005
R4099 iovss.n3098 iovss.n1167 9.0005
R4100 iovss.n3095 iovss.n1167 9.0005
R4101 iovss.n3098 iovss.n1126 9.0005
R4102 iovss.n3095 iovss.n1126 9.0005
R4103 iovss.n3098 iovss.n1170 9.0005
R4104 iovss.n3095 iovss.n1170 9.0005
R4105 iovss.n3098 iovss.n1125 9.0005
R4106 iovss.n3095 iovss.n1125 9.0005
R4107 iovss.n3098 iovss.n1173 9.0005
R4108 iovss.n3095 iovss.n1173 9.0005
R4109 iovss.n3098 iovss.n1124 9.0005
R4110 iovss.n3095 iovss.n1124 9.0005
R4111 iovss.n3098 iovss.n1175 9.0005
R4112 iovss.n3095 iovss.n1175 9.0005
R4113 iovss.n3095 iovss.n1212 9.0005
R4114 iovss.n3091 iovss.n1115 9.0005
R4115 iovss.n3095 iovss.n3091 9.0005
R4116 iovss.n3098 iovss.n1122 9.0005
R4117 iovss.n3095 iovss.n1122 9.0005
R4118 iovss.n3098 iovss.n1178 9.0005
R4119 iovss.n3095 iovss.n1178 9.0005
R4120 iovss.n3098 iovss.n1121 9.0005
R4121 iovss.n3095 iovss.n1121 9.0005
R4122 iovss.n3098 iovss.n1181 9.0005
R4123 iovss.n3095 iovss.n1181 9.0005
R4124 iovss.n3098 iovss.n1120 9.0005
R4125 iovss.n3095 iovss.n1120 9.0005
R4126 iovss.n3095 iovss.n3093 9.0005
R4127 iovss.n1210 iovss.n1115 9.0005
R4128 iovss.n3095 iovss.n1210 9.0005
R4129 iovss.n3098 iovss.n1184 9.0005
R4130 iovss.n3095 iovss.n1184 9.0005
R4131 iovss.n3098 iovss.n1119 9.0005
R4132 iovss.n3095 iovss.n1119 9.0005
R4133 iovss.n3098 iovss.n1187 9.0005
R4134 iovss.n3095 iovss.n1187 9.0005
R4135 iovss.n3098 iovss.n1118 9.0005
R4136 iovss.n3095 iovss.n1118 9.0005
R4137 iovss.n3098 iovss.n1190 9.0005
R4138 iovss.n3095 iovss.n1190 9.0005
R4139 iovss.n3098 iovss.n1117 9.0005
R4140 iovss.n3095 iovss.n1117 9.0005
R4141 iovss.n3096 iovss.n3095 9.0005
R4142 iovss.n3100 iovss.n1115 9.0005
R4143 iovss.n1103 iovss.n962 9.0005
R4144 iovss.n3109 iovss.n987 9.0005
R4145 iovss.n3109 iovss.n991 9.0005
R4146 iovss.n3109 iovss.n986 9.0005
R4147 iovss.n3109 iovss.n993 9.0005
R4148 iovss.n3109 iovss.n985 9.0005
R4149 iovss.n3109 iovss.n995 9.0005
R4150 iovss.n3109 iovss.n984 9.0005
R4151 iovss.n3109 iovss.n997 9.0005
R4152 iovss.n3109 iovss.n983 9.0005
R4153 iovss.n3109 iovss.n999 9.0005
R4154 iovss.n3109 iovss.n982 9.0005
R4155 iovss.n3109 iovss.n1001 9.0005
R4156 iovss.n3109 iovss.n981 9.0005
R4157 iovss.n3109 iovss.n1003 9.0005
R4158 iovss.n3109 iovss.n980 9.0005
R4159 iovss.n3109 iovss.n1005 9.0005
R4160 iovss.n3109 iovss.n979 9.0005
R4161 iovss.n3109 iovss.n1007 9.0005
R4162 iovss.n3109 iovss.n978 9.0005
R4163 iovss.n3109 iovss.n1009 9.0005
R4164 iovss.n3109 iovss.n977 9.0005
R4165 iovss.n3109 iovss.n1011 9.0005
R4166 iovss.n3109 iovss.n976 9.0005
R4167 iovss.n3109 iovss.n1013 9.0005
R4168 iovss.n3109 iovss.n975 9.0005
R4169 iovss.n3109 iovss.n1015 9.0005
R4170 iovss.n3109 iovss.n974 9.0005
R4171 iovss.n3109 iovss.n1017 9.0005
R4172 iovss.n3109 iovss.n973 9.0005
R4173 iovss.n3109 iovss.n1019 9.0005
R4174 iovss.n3109 iovss.n972 9.0005
R4175 iovss.n3109 iovss.n1021 9.0005
R4176 iovss.n3109 iovss.n971 9.0005
R4177 iovss.n3109 iovss.n1023 9.0005
R4178 iovss.n3109 iovss.n970 9.0005
R4179 iovss.n3109 iovss.n1025 9.0005
R4180 iovss.n3109 iovss.n969 9.0005
R4181 iovss.n3109 iovss.n1027 9.0005
R4182 iovss.n3109 iovss.n968 9.0005
R4183 iovss.n3109 iovss.n1029 9.0005
R4184 iovss.n3109 iovss.n967 9.0005
R4185 iovss.n3109 iovss.n1031 9.0005
R4186 iovss.n3109 iovss.n966 9.0005
R4187 iovss.n3109 iovss.n1033 9.0005
R4188 iovss.n3110 iovss.n3109 9.0005
R4189 iovss.n3109 iovss.n965 9.0005
R4190 iovss.n3109 iovss.n3108 9.0005
R4191 iovss.n3108 iovss.n1056 9.0005
R4192 iovss.n3108 iovss.n962 9.0005
R4193 iovss.n965 iovss.n962 9.0005
R4194 iovss.n1056 iovss.n965 9.0005
R4195 iovss.n3476 iovss.n21 9.0005
R4196 iovss.n3476 iovss.n49 9.0005
R4197 iovss.n3476 iovss.n22 9.0005
R4198 iovss.n3476 iovss.n38 9.0005
R4199 iovss.n3476 iovss.n23 9.0005
R4200 iovss.n3476 iovss.n37 9.0005
R4201 iovss.n3476 iovss.n24 9.0005
R4202 iovss.n3476 iovss.n36 9.0005
R4203 iovss.n3476 iovss.n25 9.0005
R4204 iovss.n3476 iovss.n35 9.0005
R4205 iovss.n21 iovss.n7 9.0005
R4206 iovss.n49 iovss.n7 9.0005
R4207 iovss.n22 iovss.n7 9.0005
R4208 iovss.n38 iovss.n7 9.0005
R4209 iovss.n23 iovss.n7 9.0005
R4210 iovss.n37 iovss.n7 9.0005
R4211 iovss.n24 iovss.n7 9.0005
R4212 iovss.n36 iovss.n7 9.0005
R4213 iovss.n25 iovss.n7 9.0005
R4214 iovss.n35 iovss.n7 9.0005
R4215 iovss.n31 iovss.n6 9.0005
R4216 iovss.n44 iovss.n10 9.0005
R4217 iovss.n21 iovss.n10 9.0005
R4218 iovss.n49 iovss.n10 9.0005
R4219 iovss.n22 iovss.n10 9.0005
R4220 iovss.n38 iovss.n10 9.0005
R4221 iovss.n23 iovss.n10 9.0005
R4222 iovss.n37 iovss.n10 9.0005
R4223 iovss.n24 iovss.n10 9.0005
R4224 iovss.n36 iovss.n10 9.0005
R4225 iovss.n25 iovss.n10 9.0005
R4226 iovss.n21 iovss.n11 9.0005
R4227 iovss.n49 iovss.n11 9.0005
R4228 iovss.n22 iovss.n11 9.0005
R4229 iovss.n38 iovss.n11 9.0005
R4230 iovss.n23 iovss.n11 9.0005
R4231 iovss.n37 iovss.n11 9.0005
R4232 iovss.n24 iovss.n11 9.0005
R4233 iovss.n36 iovss.n11 9.0005
R4234 iovss.n25 iovss.n11 9.0005
R4235 iovss.n35 iovss.n11 9.0005
R4236 iovss.n44 iovss.n4 9.0005
R4237 iovss.n21 iovss.n4 9.0005
R4238 iovss.n49 iovss.n4 9.0005
R4239 iovss.n22 iovss.n4 9.0005
R4240 iovss.n38 iovss.n4 9.0005
R4241 iovss.n23 iovss.n4 9.0005
R4242 iovss.n37 iovss.n4 9.0005
R4243 iovss.n24 iovss.n4 9.0005
R4244 iovss.n36 iovss.n4 9.0005
R4245 iovss.n25 iovss.n4 9.0005
R4246 iovss.n31 iovss.n12 9.0005
R4247 iovss.n21 iovss.n3 9.0005
R4248 iovss.n49 iovss.n3 9.0005
R4249 iovss.n22 iovss.n3 9.0005
R4250 iovss.n38 iovss.n3 9.0005
R4251 iovss.n23 iovss.n3 9.0005
R4252 iovss.n37 iovss.n3 9.0005
R4253 iovss.n24 iovss.n3 9.0005
R4254 iovss.n36 iovss.n3 9.0005
R4255 iovss.n25 iovss.n3 9.0005
R4256 iovss.n31 iovss.n3 9.0005
R4257 iovss.n44 iovss.n13 9.0005
R4258 iovss.n21 iovss.n13 9.0005
R4259 iovss.n49 iovss.n13 9.0005
R4260 iovss.n22 iovss.n13 9.0005
R4261 iovss.n38 iovss.n13 9.0005
R4262 iovss.n23 iovss.n13 9.0005
R4263 iovss.n37 iovss.n13 9.0005
R4264 iovss.n24 iovss.n13 9.0005
R4265 iovss.n36 iovss.n13 9.0005
R4266 iovss.n25 iovss.n13 9.0005
R4267 iovss.n21 iovss.n14 9.0005
R4268 iovss.n49 iovss.n14 9.0005
R4269 iovss.n22 iovss.n14 9.0005
R4270 iovss.n38 iovss.n14 9.0005
R4271 iovss.n23 iovss.n14 9.0005
R4272 iovss.n37 iovss.n14 9.0005
R4273 iovss.n24 iovss.n14 9.0005
R4274 iovss.n36 iovss.n14 9.0005
R4275 iovss.n25 iovss.n14 9.0005
R4276 iovss.n35 iovss.n14 9.0005
R4277 iovss.n44 iovss.n1 9.0005
R4278 iovss.n21 iovss.n1 9.0005
R4279 iovss.n49 iovss.n1 9.0005
R4280 iovss.n22 iovss.n1 9.0005
R4281 iovss.n38 iovss.n1 9.0005
R4282 iovss.n23 iovss.n1 9.0005
R4283 iovss.n37 iovss.n1 9.0005
R4284 iovss.n24 iovss.n1 9.0005
R4285 iovss.n36 iovss.n1 9.0005
R4286 iovss.n25 iovss.n1 9.0005
R4287 iovss.n35 iovss.n1 9.0005
R4288 iovss.n35 iovss.n2 9.0005
R4289 iovss.n25 iovss.n2 9.0005
R4290 iovss.n36 iovss.n2 9.0005
R4291 iovss.n24 iovss.n2 9.0005
R4292 iovss.n37 iovss.n2 9.0005
R4293 iovss.n23 iovss.n2 9.0005
R4294 iovss.n38 iovss.n2 9.0005
R4295 iovss.n22 iovss.n2 9.0005
R4296 iovss.n49 iovss.n2 9.0005
R4297 iovss.n21 iovss.n2 9.0005
R4298 iovss.n25 iovss.n12 9.0005
R4299 iovss.n36 iovss.n12 9.0005
R4300 iovss.n24 iovss.n12 9.0005
R4301 iovss.n37 iovss.n12 9.0005
R4302 iovss.n23 iovss.n12 9.0005
R4303 iovss.n38 iovss.n12 9.0005
R4304 iovss.n22 iovss.n12 9.0005
R4305 iovss.n49 iovss.n12 9.0005
R4306 iovss.n21 iovss.n12 9.0005
R4307 iovss.n35 iovss.n5 9.0005
R4308 iovss.n25 iovss.n5 9.0005
R4309 iovss.n36 iovss.n5 9.0005
R4310 iovss.n24 iovss.n5 9.0005
R4311 iovss.n37 iovss.n5 9.0005
R4312 iovss.n23 iovss.n5 9.0005
R4313 iovss.n38 iovss.n5 9.0005
R4314 iovss.n22 iovss.n5 9.0005
R4315 iovss.n49 iovss.n5 9.0005
R4316 iovss.n21 iovss.n5 9.0005
R4317 iovss.n25 iovss.n6 9.0005
R4318 iovss.n36 iovss.n6 9.0005
R4319 iovss.n24 iovss.n6 9.0005
R4320 iovss.n37 iovss.n6 9.0005
R4321 iovss.n23 iovss.n6 9.0005
R4322 iovss.n38 iovss.n6 9.0005
R4323 iovss.n22 iovss.n6 9.0005
R4324 iovss.n49 iovss.n6 9.0005
R4325 iovss.n21 iovss.n6 9.0005
R4326 iovss.n35 iovss.n9 9.0005
R4327 iovss.n25 iovss.n9 9.0005
R4328 iovss.n36 iovss.n9 9.0005
R4329 iovss.n24 iovss.n9 9.0005
R4330 iovss.n37 iovss.n9 9.0005
R4331 iovss.n23 iovss.n9 9.0005
R4332 iovss.n38 iovss.n9 9.0005
R4333 iovss.n22 iovss.n9 9.0005
R4334 iovss.n49 iovss.n9 9.0005
R4335 iovss.n21 iovss.n9 9.0005
R4336 iovss.n35 iovss.n8 9.0005
R4337 iovss.n25 iovss.n8 9.0005
R4338 iovss.n36 iovss.n8 9.0005
R4339 iovss.n24 iovss.n8 9.0005
R4340 iovss.n37 iovss.n8 9.0005
R4341 iovss.n23 iovss.n8 9.0005
R4342 iovss.n38 iovss.n8 9.0005
R4343 iovss.n22 iovss.n8 9.0005
R4344 iovss.n49 iovss.n8 9.0005
R4345 iovss.n21 iovss.n8 9.0005
R4346 iovss.n3479 iovss.n31 9.0005
R4347 iovss.n3479 iovss.n35 9.0005
R4348 iovss.n3479 iovss.n25 9.0005
R4349 iovss.n3479 iovss.n36 9.0005
R4350 iovss.n3479 iovss.n24 9.0005
R4351 iovss.n3479 iovss.n37 9.0005
R4352 iovss.n3479 iovss.n23 9.0005
R4353 iovss.n3479 iovss.n38 9.0005
R4354 iovss.n3479 iovss.n22 9.0005
R4355 iovss.n3479 iovss.n49 9.0005
R4356 iovss.n3479 iovss.n21 9.0005
R4357 iovss.n3254 iovss.n530 9.0005
R4358 iovss.n537 iovss.n498 9.0005
R4359 iovss.n538 iovss.n498 9.0005
R4360 iovss.n536 iovss.n498 9.0005
R4361 iovss.n541 iovss.n498 9.0005
R4362 iovss.n534 iovss.n498 9.0005
R4363 iovss.n544 iovss.n498 9.0005
R4364 iovss.n532 iovss.n498 9.0005
R4365 iovss.n547 iovss.n498 9.0005
R4366 iovss.n528 iovss.n498 9.0005
R4367 iovss.n552 iovss.n498 9.0005
R4368 iovss.n526 iovss.n498 9.0005
R4369 iovss.n555 iovss.n498 9.0005
R4370 iovss.n524 iovss.n498 9.0005
R4371 iovss.n609 iovss.n498 9.0005
R4372 iovss.n522 iovss.n498 9.0005
R4373 iovss.n613 iovss.n498 9.0005
R4374 iovss.n498 iovss.n489 9.0005
R4375 iovss.n3259 iovss.n498 9.0005
R4376 iovss.n537 iovss.n496 9.0005
R4377 iovss.n538 iovss.n496 9.0005
R4378 iovss.n536 iovss.n496 9.0005
R4379 iovss.n540 iovss.n496 9.0005
R4380 iovss.n535 iovss.n496 9.0005
R4381 iovss.n541 iovss.n496 9.0005
R4382 iovss.n534 iovss.n496 9.0005
R4383 iovss.n543 iovss.n496 9.0005
R4384 iovss.n533 iovss.n496 9.0005
R4385 iovss.n544 iovss.n496 9.0005
R4386 iovss.n532 iovss.n496 9.0005
R4387 iovss.n546 iovss.n496 9.0005
R4388 iovss.n531 iovss.n496 9.0005
R4389 iovss.n547 iovss.n496 9.0005
R4390 iovss.n530 iovss.n496 9.0005
R4391 iovss.n549 iovss.n496 9.0005
R4392 iovss.n529 iovss.n496 9.0005
R4393 iovss.n551 iovss.n496 9.0005
R4394 iovss.n528 iovss.n496 9.0005
R4395 iovss.n552 iovss.n496 9.0005
R4396 iovss.n527 iovss.n496 9.0005
R4397 iovss.n554 iovss.n496 9.0005
R4398 iovss.n526 iovss.n496 9.0005
R4399 iovss.n555 iovss.n496 9.0005
R4400 iovss.n525 iovss.n496 9.0005
R4401 iovss.n557 iovss.n496 9.0005
R4402 iovss.n524 iovss.n496 9.0005
R4403 iovss.n609 iovss.n496 9.0005
R4404 iovss.n523 iovss.n496 9.0005
R4405 iovss.n611 iovss.n496 9.0005
R4406 iovss.n522 iovss.n496 9.0005
R4407 iovss.n613 iovss.n496 9.0005
R4408 iovss.n521 iovss.n496 9.0005
R4409 iovss.n3257 iovss.n496 9.0005
R4410 iovss.n3259 iovss.n496 9.0005
R4411 iovss.n614 iovss.n496 9.0005
R4412 iovss.n537 iovss.n500 9.0005
R4413 iovss.n538 iovss.n500 9.0005
R4414 iovss.n536 iovss.n500 9.0005
R4415 iovss.n540 iovss.n500 9.0005
R4416 iovss.n535 iovss.n500 9.0005
R4417 iovss.n541 iovss.n500 9.0005
R4418 iovss.n534 iovss.n500 9.0005
R4419 iovss.n543 iovss.n500 9.0005
R4420 iovss.n533 iovss.n500 9.0005
R4421 iovss.n544 iovss.n500 9.0005
R4422 iovss.n532 iovss.n500 9.0005
R4423 iovss.n546 iovss.n500 9.0005
R4424 iovss.n531 iovss.n500 9.0005
R4425 iovss.n547 iovss.n500 9.0005
R4426 iovss.n530 iovss.n500 9.0005
R4427 iovss.n549 iovss.n500 9.0005
R4428 iovss.n529 iovss.n500 9.0005
R4429 iovss.n551 iovss.n500 9.0005
R4430 iovss.n528 iovss.n500 9.0005
R4431 iovss.n552 iovss.n500 9.0005
R4432 iovss.n527 iovss.n500 9.0005
R4433 iovss.n554 iovss.n500 9.0005
R4434 iovss.n526 iovss.n500 9.0005
R4435 iovss.n555 iovss.n500 9.0005
R4436 iovss.n525 iovss.n500 9.0005
R4437 iovss.n557 iovss.n500 9.0005
R4438 iovss.n524 iovss.n500 9.0005
R4439 iovss.n609 iovss.n500 9.0005
R4440 iovss.n523 iovss.n500 9.0005
R4441 iovss.n611 iovss.n500 9.0005
R4442 iovss.n522 iovss.n500 9.0005
R4443 iovss.n613 iovss.n500 9.0005
R4444 iovss.n521 iovss.n500 9.0005
R4445 iovss.n3257 iovss.n500 9.0005
R4446 iovss.n3259 iovss.n500 9.0005
R4447 iovss.n614 iovss.n500 9.0005
R4448 iovss.n537 iovss.n495 9.0005
R4449 iovss.n538 iovss.n495 9.0005
R4450 iovss.n536 iovss.n495 9.0005
R4451 iovss.n540 iovss.n495 9.0005
R4452 iovss.n535 iovss.n495 9.0005
R4453 iovss.n541 iovss.n495 9.0005
R4454 iovss.n534 iovss.n495 9.0005
R4455 iovss.n543 iovss.n495 9.0005
R4456 iovss.n533 iovss.n495 9.0005
R4457 iovss.n544 iovss.n495 9.0005
R4458 iovss.n532 iovss.n495 9.0005
R4459 iovss.n546 iovss.n495 9.0005
R4460 iovss.n531 iovss.n495 9.0005
R4461 iovss.n547 iovss.n495 9.0005
R4462 iovss.n530 iovss.n495 9.0005
R4463 iovss.n549 iovss.n495 9.0005
R4464 iovss.n529 iovss.n495 9.0005
R4465 iovss.n551 iovss.n495 9.0005
R4466 iovss.n528 iovss.n495 9.0005
R4467 iovss.n552 iovss.n495 9.0005
R4468 iovss.n527 iovss.n495 9.0005
R4469 iovss.n554 iovss.n495 9.0005
R4470 iovss.n526 iovss.n495 9.0005
R4471 iovss.n555 iovss.n495 9.0005
R4472 iovss.n525 iovss.n495 9.0005
R4473 iovss.n557 iovss.n495 9.0005
R4474 iovss.n524 iovss.n495 9.0005
R4475 iovss.n609 iovss.n495 9.0005
R4476 iovss.n523 iovss.n495 9.0005
R4477 iovss.n611 iovss.n495 9.0005
R4478 iovss.n522 iovss.n495 9.0005
R4479 iovss.n613 iovss.n495 9.0005
R4480 iovss.n521 iovss.n495 9.0005
R4481 iovss.n3257 iovss.n495 9.0005
R4482 iovss.n3259 iovss.n495 9.0005
R4483 iovss.n614 iovss.n495 9.0005
R4484 iovss.n537 iovss.n502 9.0005
R4485 iovss.n538 iovss.n502 9.0005
R4486 iovss.n536 iovss.n502 9.0005
R4487 iovss.n540 iovss.n502 9.0005
R4488 iovss.n535 iovss.n502 9.0005
R4489 iovss.n541 iovss.n502 9.0005
R4490 iovss.n534 iovss.n502 9.0005
R4491 iovss.n543 iovss.n502 9.0005
R4492 iovss.n533 iovss.n502 9.0005
R4493 iovss.n544 iovss.n502 9.0005
R4494 iovss.n532 iovss.n502 9.0005
R4495 iovss.n546 iovss.n502 9.0005
R4496 iovss.n531 iovss.n502 9.0005
R4497 iovss.n547 iovss.n502 9.0005
R4498 iovss.n530 iovss.n502 9.0005
R4499 iovss.n549 iovss.n502 9.0005
R4500 iovss.n529 iovss.n502 9.0005
R4501 iovss.n551 iovss.n502 9.0005
R4502 iovss.n528 iovss.n502 9.0005
R4503 iovss.n552 iovss.n502 9.0005
R4504 iovss.n527 iovss.n502 9.0005
R4505 iovss.n554 iovss.n502 9.0005
R4506 iovss.n526 iovss.n502 9.0005
R4507 iovss.n555 iovss.n502 9.0005
R4508 iovss.n525 iovss.n502 9.0005
R4509 iovss.n557 iovss.n502 9.0005
R4510 iovss.n524 iovss.n502 9.0005
R4511 iovss.n609 iovss.n502 9.0005
R4512 iovss.n523 iovss.n502 9.0005
R4513 iovss.n611 iovss.n502 9.0005
R4514 iovss.n522 iovss.n502 9.0005
R4515 iovss.n613 iovss.n502 9.0005
R4516 iovss.n521 iovss.n502 9.0005
R4517 iovss.n3257 iovss.n502 9.0005
R4518 iovss.n3259 iovss.n502 9.0005
R4519 iovss.n614 iovss.n502 9.0005
R4520 iovss.n537 iovss.n494 9.0005
R4521 iovss.n538 iovss.n494 9.0005
R4522 iovss.n536 iovss.n494 9.0005
R4523 iovss.n540 iovss.n494 9.0005
R4524 iovss.n535 iovss.n494 9.0005
R4525 iovss.n541 iovss.n494 9.0005
R4526 iovss.n534 iovss.n494 9.0005
R4527 iovss.n543 iovss.n494 9.0005
R4528 iovss.n533 iovss.n494 9.0005
R4529 iovss.n544 iovss.n494 9.0005
R4530 iovss.n532 iovss.n494 9.0005
R4531 iovss.n546 iovss.n494 9.0005
R4532 iovss.n531 iovss.n494 9.0005
R4533 iovss.n547 iovss.n494 9.0005
R4534 iovss.n530 iovss.n494 9.0005
R4535 iovss.n549 iovss.n494 9.0005
R4536 iovss.n529 iovss.n494 9.0005
R4537 iovss.n551 iovss.n494 9.0005
R4538 iovss.n528 iovss.n494 9.0005
R4539 iovss.n552 iovss.n494 9.0005
R4540 iovss.n527 iovss.n494 9.0005
R4541 iovss.n554 iovss.n494 9.0005
R4542 iovss.n526 iovss.n494 9.0005
R4543 iovss.n555 iovss.n494 9.0005
R4544 iovss.n525 iovss.n494 9.0005
R4545 iovss.n557 iovss.n494 9.0005
R4546 iovss.n524 iovss.n494 9.0005
R4547 iovss.n609 iovss.n494 9.0005
R4548 iovss.n523 iovss.n494 9.0005
R4549 iovss.n611 iovss.n494 9.0005
R4550 iovss.n522 iovss.n494 9.0005
R4551 iovss.n613 iovss.n494 9.0005
R4552 iovss.n521 iovss.n494 9.0005
R4553 iovss.n3257 iovss.n494 9.0005
R4554 iovss.n3259 iovss.n494 9.0005
R4555 iovss.n614 iovss.n494 9.0005
R4556 iovss.n537 iovss.n504 9.0005
R4557 iovss.n538 iovss.n504 9.0005
R4558 iovss.n536 iovss.n504 9.0005
R4559 iovss.n540 iovss.n504 9.0005
R4560 iovss.n535 iovss.n504 9.0005
R4561 iovss.n541 iovss.n504 9.0005
R4562 iovss.n534 iovss.n504 9.0005
R4563 iovss.n543 iovss.n504 9.0005
R4564 iovss.n533 iovss.n504 9.0005
R4565 iovss.n544 iovss.n504 9.0005
R4566 iovss.n532 iovss.n504 9.0005
R4567 iovss.n546 iovss.n504 9.0005
R4568 iovss.n531 iovss.n504 9.0005
R4569 iovss.n547 iovss.n504 9.0005
R4570 iovss.n530 iovss.n504 9.0005
R4571 iovss.n549 iovss.n504 9.0005
R4572 iovss.n529 iovss.n504 9.0005
R4573 iovss.n551 iovss.n504 9.0005
R4574 iovss.n528 iovss.n504 9.0005
R4575 iovss.n552 iovss.n504 9.0005
R4576 iovss.n527 iovss.n504 9.0005
R4577 iovss.n554 iovss.n504 9.0005
R4578 iovss.n526 iovss.n504 9.0005
R4579 iovss.n555 iovss.n504 9.0005
R4580 iovss.n525 iovss.n504 9.0005
R4581 iovss.n557 iovss.n504 9.0005
R4582 iovss.n524 iovss.n504 9.0005
R4583 iovss.n609 iovss.n504 9.0005
R4584 iovss.n523 iovss.n504 9.0005
R4585 iovss.n611 iovss.n504 9.0005
R4586 iovss.n522 iovss.n504 9.0005
R4587 iovss.n613 iovss.n504 9.0005
R4588 iovss.n521 iovss.n504 9.0005
R4589 iovss.n3257 iovss.n504 9.0005
R4590 iovss.n3259 iovss.n504 9.0005
R4591 iovss.n614 iovss.n504 9.0005
R4592 iovss.n537 iovss.n493 9.0005
R4593 iovss.n538 iovss.n493 9.0005
R4594 iovss.n536 iovss.n493 9.0005
R4595 iovss.n540 iovss.n493 9.0005
R4596 iovss.n535 iovss.n493 9.0005
R4597 iovss.n541 iovss.n493 9.0005
R4598 iovss.n534 iovss.n493 9.0005
R4599 iovss.n543 iovss.n493 9.0005
R4600 iovss.n533 iovss.n493 9.0005
R4601 iovss.n544 iovss.n493 9.0005
R4602 iovss.n532 iovss.n493 9.0005
R4603 iovss.n546 iovss.n493 9.0005
R4604 iovss.n531 iovss.n493 9.0005
R4605 iovss.n547 iovss.n493 9.0005
R4606 iovss.n530 iovss.n493 9.0005
R4607 iovss.n549 iovss.n493 9.0005
R4608 iovss.n529 iovss.n493 9.0005
R4609 iovss.n551 iovss.n493 9.0005
R4610 iovss.n528 iovss.n493 9.0005
R4611 iovss.n552 iovss.n493 9.0005
R4612 iovss.n527 iovss.n493 9.0005
R4613 iovss.n554 iovss.n493 9.0005
R4614 iovss.n526 iovss.n493 9.0005
R4615 iovss.n555 iovss.n493 9.0005
R4616 iovss.n525 iovss.n493 9.0005
R4617 iovss.n557 iovss.n493 9.0005
R4618 iovss.n524 iovss.n493 9.0005
R4619 iovss.n609 iovss.n493 9.0005
R4620 iovss.n523 iovss.n493 9.0005
R4621 iovss.n611 iovss.n493 9.0005
R4622 iovss.n522 iovss.n493 9.0005
R4623 iovss.n613 iovss.n493 9.0005
R4624 iovss.n521 iovss.n493 9.0005
R4625 iovss.n3257 iovss.n493 9.0005
R4626 iovss.n3259 iovss.n493 9.0005
R4627 iovss.n614 iovss.n493 9.0005
R4628 iovss.n537 iovss.n506 9.0005
R4629 iovss.n538 iovss.n506 9.0005
R4630 iovss.n536 iovss.n506 9.0005
R4631 iovss.n540 iovss.n506 9.0005
R4632 iovss.n535 iovss.n506 9.0005
R4633 iovss.n541 iovss.n506 9.0005
R4634 iovss.n534 iovss.n506 9.0005
R4635 iovss.n543 iovss.n506 9.0005
R4636 iovss.n533 iovss.n506 9.0005
R4637 iovss.n544 iovss.n506 9.0005
R4638 iovss.n532 iovss.n506 9.0005
R4639 iovss.n546 iovss.n506 9.0005
R4640 iovss.n531 iovss.n506 9.0005
R4641 iovss.n547 iovss.n506 9.0005
R4642 iovss.n530 iovss.n506 9.0005
R4643 iovss.n549 iovss.n506 9.0005
R4644 iovss.n529 iovss.n506 9.0005
R4645 iovss.n551 iovss.n506 9.0005
R4646 iovss.n528 iovss.n506 9.0005
R4647 iovss.n552 iovss.n506 9.0005
R4648 iovss.n527 iovss.n506 9.0005
R4649 iovss.n554 iovss.n506 9.0005
R4650 iovss.n526 iovss.n506 9.0005
R4651 iovss.n555 iovss.n506 9.0005
R4652 iovss.n525 iovss.n506 9.0005
R4653 iovss.n557 iovss.n506 9.0005
R4654 iovss.n524 iovss.n506 9.0005
R4655 iovss.n609 iovss.n506 9.0005
R4656 iovss.n523 iovss.n506 9.0005
R4657 iovss.n611 iovss.n506 9.0005
R4658 iovss.n522 iovss.n506 9.0005
R4659 iovss.n613 iovss.n506 9.0005
R4660 iovss.n521 iovss.n506 9.0005
R4661 iovss.n3257 iovss.n506 9.0005
R4662 iovss.n3259 iovss.n506 9.0005
R4663 iovss.n614 iovss.n506 9.0005
R4664 iovss.n537 iovss.n492 9.0005
R4665 iovss.n538 iovss.n492 9.0005
R4666 iovss.n536 iovss.n492 9.0005
R4667 iovss.n540 iovss.n492 9.0005
R4668 iovss.n535 iovss.n492 9.0005
R4669 iovss.n541 iovss.n492 9.0005
R4670 iovss.n534 iovss.n492 9.0005
R4671 iovss.n543 iovss.n492 9.0005
R4672 iovss.n533 iovss.n492 9.0005
R4673 iovss.n544 iovss.n492 9.0005
R4674 iovss.n532 iovss.n492 9.0005
R4675 iovss.n546 iovss.n492 9.0005
R4676 iovss.n531 iovss.n492 9.0005
R4677 iovss.n547 iovss.n492 9.0005
R4678 iovss.n530 iovss.n492 9.0005
R4679 iovss.n549 iovss.n492 9.0005
R4680 iovss.n529 iovss.n492 9.0005
R4681 iovss.n551 iovss.n492 9.0005
R4682 iovss.n528 iovss.n492 9.0005
R4683 iovss.n552 iovss.n492 9.0005
R4684 iovss.n527 iovss.n492 9.0005
R4685 iovss.n554 iovss.n492 9.0005
R4686 iovss.n526 iovss.n492 9.0005
R4687 iovss.n555 iovss.n492 9.0005
R4688 iovss.n525 iovss.n492 9.0005
R4689 iovss.n557 iovss.n492 9.0005
R4690 iovss.n524 iovss.n492 9.0005
R4691 iovss.n609 iovss.n492 9.0005
R4692 iovss.n523 iovss.n492 9.0005
R4693 iovss.n611 iovss.n492 9.0005
R4694 iovss.n522 iovss.n492 9.0005
R4695 iovss.n613 iovss.n492 9.0005
R4696 iovss.n521 iovss.n492 9.0005
R4697 iovss.n3257 iovss.n492 9.0005
R4698 iovss.n3259 iovss.n492 9.0005
R4699 iovss.n614 iovss.n492 9.0005
R4700 iovss.n537 iovss.n508 9.0005
R4701 iovss.n538 iovss.n508 9.0005
R4702 iovss.n536 iovss.n508 9.0005
R4703 iovss.n540 iovss.n508 9.0005
R4704 iovss.n535 iovss.n508 9.0005
R4705 iovss.n541 iovss.n508 9.0005
R4706 iovss.n534 iovss.n508 9.0005
R4707 iovss.n543 iovss.n508 9.0005
R4708 iovss.n533 iovss.n508 9.0005
R4709 iovss.n544 iovss.n508 9.0005
R4710 iovss.n532 iovss.n508 9.0005
R4711 iovss.n546 iovss.n508 9.0005
R4712 iovss.n531 iovss.n508 9.0005
R4713 iovss.n547 iovss.n508 9.0005
R4714 iovss.n530 iovss.n508 9.0005
R4715 iovss.n549 iovss.n508 9.0005
R4716 iovss.n529 iovss.n508 9.0005
R4717 iovss.n551 iovss.n508 9.0005
R4718 iovss.n528 iovss.n508 9.0005
R4719 iovss.n552 iovss.n508 9.0005
R4720 iovss.n527 iovss.n508 9.0005
R4721 iovss.n554 iovss.n508 9.0005
R4722 iovss.n526 iovss.n508 9.0005
R4723 iovss.n555 iovss.n508 9.0005
R4724 iovss.n525 iovss.n508 9.0005
R4725 iovss.n557 iovss.n508 9.0005
R4726 iovss.n524 iovss.n508 9.0005
R4727 iovss.n609 iovss.n508 9.0005
R4728 iovss.n523 iovss.n508 9.0005
R4729 iovss.n611 iovss.n508 9.0005
R4730 iovss.n522 iovss.n508 9.0005
R4731 iovss.n613 iovss.n508 9.0005
R4732 iovss.n521 iovss.n508 9.0005
R4733 iovss.n3257 iovss.n508 9.0005
R4734 iovss.n3259 iovss.n508 9.0005
R4735 iovss.n614 iovss.n508 9.0005
R4736 iovss.n537 iovss.n491 9.0005
R4737 iovss.n538 iovss.n491 9.0005
R4738 iovss.n536 iovss.n491 9.0005
R4739 iovss.n540 iovss.n491 9.0005
R4740 iovss.n535 iovss.n491 9.0005
R4741 iovss.n541 iovss.n491 9.0005
R4742 iovss.n534 iovss.n491 9.0005
R4743 iovss.n543 iovss.n491 9.0005
R4744 iovss.n533 iovss.n491 9.0005
R4745 iovss.n544 iovss.n491 9.0005
R4746 iovss.n532 iovss.n491 9.0005
R4747 iovss.n546 iovss.n491 9.0005
R4748 iovss.n531 iovss.n491 9.0005
R4749 iovss.n547 iovss.n491 9.0005
R4750 iovss.n530 iovss.n491 9.0005
R4751 iovss.n549 iovss.n491 9.0005
R4752 iovss.n529 iovss.n491 9.0005
R4753 iovss.n551 iovss.n491 9.0005
R4754 iovss.n528 iovss.n491 9.0005
R4755 iovss.n552 iovss.n491 9.0005
R4756 iovss.n527 iovss.n491 9.0005
R4757 iovss.n554 iovss.n491 9.0005
R4758 iovss.n526 iovss.n491 9.0005
R4759 iovss.n555 iovss.n491 9.0005
R4760 iovss.n525 iovss.n491 9.0005
R4761 iovss.n557 iovss.n491 9.0005
R4762 iovss.n524 iovss.n491 9.0005
R4763 iovss.n609 iovss.n491 9.0005
R4764 iovss.n523 iovss.n491 9.0005
R4765 iovss.n611 iovss.n491 9.0005
R4766 iovss.n522 iovss.n491 9.0005
R4767 iovss.n613 iovss.n491 9.0005
R4768 iovss.n521 iovss.n491 9.0005
R4769 iovss.n3257 iovss.n491 9.0005
R4770 iovss.n3259 iovss.n491 9.0005
R4771 iovss.n614 iovss.n491 9.0005
R4772 iovss.n537 iovss.n510 9.0005
R4773 iovss.n538 iovss.n510 9.0005
R4774 iovss.n536 iovss.n510 9.0005
R4775 iovss.n540 iovss.n510 9.0005
R4776 iovss.n535 iovss.n510 9.0005
R4777 iovss.n541 iovss.n510 9.0005
R4778 iovss.n534 iovss.n510 9.0005
R4779 iovss.n543 iovss.n510 9.0005
R4780 iovss.n533 iovss.n510 9.0005
R4781 iovss.n544 iovss.n510 9.0005
R4782 iovss.n532 iovss.n510 9.0005
R4783 iovss.n546 iovss.n510 9.0005
R4784 iovss.n531 iovss.n510 9.0005
R4785 iovss.n547 iovss.n510 9.0005
R4786 iovss.n530 iovss.n510 9.0005
R4787 iovss.n549 iovss.n510 9.0005
R4788 iovss.n529 iovss.n510 9.0005
R4789 iovss.n551 iovss.n510 9.0005
R4790 iovss.n528 iovss.n510 9.0005
R4791 iovss.n552 iovss.n510 9.0005
R4792 iovss.n527 iovss.n510 9.0005
R4793 iovss.n554 iovss.n510 9.0005
R4794 iovss.n526 iovss.n510 9.0005
R4795 iovss.n555 iovss.n510 9.0005
R4796 iovss.n525 iovss.n510 9.0005
R4797 iovss.n557 iovss.n510 9.0005
R4798 iovss.n524 iovss.n510 9.0005
R4799 iovss.n609 iovss.n510 9.0005
R4800 iovss.n523 iovss.n510 9.0005
R4801 iovss.n611 iovss.n510 9.0005
R4802 iovss.n522 iovss.n510 9.0005
R4803 iovss.n613 iovss.n510 9.0005
R4804 iovss.n521 iovss.n510 9.0005
R4805 iovss.n3257 iovss.n510 9.0005
R4806 iovss.n3259 iovss.n510 9.0005
R4807 iovss.n614 iovss.n510 9.0005
R4808 iovss.n537 iovss.n490 9.0005
R4809 iovss.n538 iovss.n490 9.0005
R4810 iovss.n536 iovss.n490 9.0005
R4811 iovss.n540 iovss.n490 9.0005
R4812 iovss.n535 iovss.n490 9.0005
R4813 iovss.n541 iovss.n490 9.0005
R4814 iovss.n534 iovss.n490 9.0005
R4815 iovss.n543 iovss.n490 9.0005
R4816 iovss.n533 iovss.n490 9.0005
R4817 iovss.n544 iovss.n490 9.0005
R4818 iovss.n532 iovss.n490 9.0005
R4819 iovss.n546 iovss.n490 9.0005
R4820 iovss.n531 iovss.n490 9.0005
R4821 iovss.n547 iovss.n490 9.0005
R4822 iovss.n530 iovss.n490 9.0005
R4823 iovss.n549 iovss.n490 9.0005
R4824 iovss.n529 iovss.n490 9.0005
R4825 iovss.n551 iovss.n490 9.0005
R4826 iovss.n528 iovss.n490 9.0005
R4827 iovss.n552 iovss.n490 9.0005
R4828 iovss.n527 iovss.n490 9.0005
R4829 iovss.n554 iovss.n490 9.0005
R4830 iovss.n526 iovss.n490 9.0005
R4831 iovss.n555 iovss.n490 9.0005
R4832 iovss.n525 iovss.n490 9.0005
R4833 iovss.n557 iovss.n490 9.0005
R4834 iovss.n524 iovss.n490 9.0005
R4835 iovss.n609 iovss.n490 9.0005
R4836 iovss.n523 iovss.n490 9.0005
R4837 iovss.n611 iovss.n490 9.0005
R4838 iovss.n522 iovss.n490 9.0005
R4839 iovss.n613 iovss.n490 9.0005
R4840 iovss.n521 iovss.n490 9.0005
R4841 iovss.n3257 iovss.n490 9.0005
R4842 iovss.n3259 iovss.n490 9.0005
R4843 iovss.n614 iovss.n490 9.0005
R4844 iovss.n3258 iovss.n537 9.0005
R4845 iovss.n3258 iovss.n538 9.0005
R4846 iovss.n3258 iovss.n536 9.0005
R4847 iovss.n3258 iovss.n540 9.0005
R4848 iovss.n3258 iovss.n535 9.0005
R4849 iovss.n3258 iovss.n541 9.0005
R4850 iovss.n3258 iovss.n534 9.0005
R4851 iovss.n3258 iovss.n543 9.0005
R4852 iovss.n3258 iovss.n533 9.0005
R4853 iovss.n3258 iovss.n544 9.0005
R4854 iovss.n3258 iovss.n532 9.0005
R4855 iovss.n3258 iovss.n546 9.0005
R4856 iovss.n3258 iovss.n531 9.0005
R4857 iovss.n3258 iovss.n547 9.0005
R4858 iovss.n3258 iovss.n530 9.0005
R4859 iovss.n3258 iovss.n549 9.0005
R4860 iovss.n3258 iovss.n529 9.0005
R4861 iovss.n3258 iovss.n551 9.0005
R4862 iovss.n3258 iovss.n528 9.0005
R4863 iovss.n3258 iovss.n552 9.0005
R4864 iovss.n3258 iovss.n527 9.0005
R4865 iovss.n3258 iovss.n554 9.0005
R4866 iovss.n3258 iovss.n526 9.0005
R4867 iovss.n3258 iovss.n555 9.0005
R4868 iovss.n3258 iovss.n525 9.0005
R4869 iovss.n3258 iovss.n557 9.0005
R4870 iovss.n3258 iovss.n524 9.0005
R4871 iovss.n3258 iovss.n609 9.0005
R4872 iovss.n3258 iovss.n523 9.0005
R4873 iovss.n3258 iovss.n611 9.0005
R4874 iovss.n3258 iovss.n522 9.0005
R4875 iovss.n3258 iovss.n613 9.0005
R4876 iovss.n3258 iovss.n521 9.0005
R4877 iovss.n3258 iovss.n3257 9.0005
R4878 iovss.n3259 iovss.n3258 9.0005
R4879 iovss.n3344 iovss.n3343 9.0005
R4880 iovss.n3344 iovss.n373 9.0005
R4881 iovss.n3344 iovss.n362 9.0005
R4882 iovss.n3343 iovss.n389 9.0005
R4883 iovss.n429 iovss.n389 9.0005
R4884 iovss.n427 iovss.n389 9.0005
R4885 iovss.n432 iovss.n389 9.0005
R4886 iovss.n425 iovss.n389 9.0005
R4887 iovss.n435 iovss.n389 9.0005
R4888 iovss.n423 iovss.n389 9.0005
R4889 iovss.n440 iovss.n389 9.0005
R4890 iovss.n419 iovss.n389 9.0005
R4891 iovss.n443 iovss.n389 9.0005
R4892 iovss.n417 iovss.n389 9.0005
R4893 iovss.n446 iovss.n389 9.0005
R4894 iovss.n415 iovss.n389 9.0005
R4895 iovss.n449 iovss.n389 9.0005
R4896 iovss.n413 iovss.n389 9.0005
R4897 iovss.n3339 iovss.n389 9.0005
R4898 iovss.n3343 iovss.n387 9.0005
R4899 iovss.n429 iovss.n387 9.0005
R4900 iovss.n428 iovss.n387 9.0005
R4901 iovss.n431 iovss.n387 9.0005
R4902 iovss.n427 iovss.n387 9.0005
R4903 iovss.n432 iovss.n387 9.0005
R4904 iovss.n426 iovss.n387 9.0005
R4905 iovss.n434 iovss.n387 9.0005
R4906 iovss.n425 iovss.n387 9.0005
R4907 iovss.n435 iovss.n387 9.0005
R4908 iovss.n424 iovss.n387 9.0005
R4909 iovss.n437 iovss.n387 9.0005
R4910 iovss.n423 iovss.n387 9.0005
R4911 iovss.n387 iovss.n373 9.0005
R4912 iovss.n422 iovss.n387 9.0005
R4913 iovss.n439 iovss.n387 9.0005
R4914 iovss.n420 iovss.n387 9.0005
R4915 iovss.n440 iovss.n387 9.0005
R4916 iovss.n419 iovss.n387 9.0005
R4917 iovss.n442 iovss.n387 9.0005
R4918 iovss.n418 iovss.n387 9.0005
R4919 iovss.n443 iovss.n387 9.0005
R4920 iovss.n417 iovss.n387 9.0005
R4921 iovss.n445 iovss.n387 9.0005
R4922 iovss.n416 iovss.n387 9.0005
R4923 iovss.n446 iovss.n387 9.0005
R4924 iovss.n415 iovss.n387 9.0005
R4925 iovss.n448 iovss.n387 9.0005
R4926 iovss.n414 iovss.n387 9.0005
R4927 iovss.n449 iovss.n387 9.0005
R4928 iovss.n413 iovss.n387 9.0005
R4929 iovss.n451 iovss.n387 9.0005
R4930 iovss.n412 iovss.n387 9.0005
R4931 iovss.n3339 iovss.n387 9.0005
R4932 iovss.n3341 iovss.n387 9.0005
R4933 iovss.n3333 iovss.n387 9.0005
R4934 iovss.n3343 iovss.n391 9.0005
R4935 iovss.n429 iovss.n391 9.0005
R4936 iovss.n428 iovss.n391 9.0005
R4937 iovss.n431 iovss.n391 9.0005
R4938 iovss.n427 iovss.n391 9.0005
R4939 iovss.n432 iovss.n391 9.0005
R4940 iovss.n426 iovss.n391 9.0005
R4941 iovss.n434 iovss.n391 9.0005
R4942 iovss.n425 iovss.n391 9.0005
R4943 iovss.n435 iovss.n391 9.0005
R4944 iovss.n424 iovss.n391 9.0005
R4945 iovss.n437 iovss.n391 9.0005
R4946 iovss.n423 iovss.n391 9.0005
R4947 iovss.n391 iovss.n373 9.0005
R4948 iovss.n422 iovss.n391 9.0005
R4949 iovss.n439 iovss.n391 9.0005
R4950 iovss.n420 iovss.n391 9.0005
R4951 iovss.n440 iovss.n391 9.0005
R4952 iovss.n419 iovss.n391 9.0005
R4953 iovss.n442 iovss.n391 9.0005
R4954 iovss.n418 iovss.n391 9.0005
R4955 iovss.n443 iovss.n391 9.0005
R4956 iovss.n417 iovss.n391 9.0005
R4957 iovss.n445 iovss.n391 9.0005
R4958 iovss.n416 iovss.n391 9.0005
R4959 iovss.n446 iovss.n391 9.0005
R4960 iovss.n415 iovss.n391 9.0005
R4961 iovss.n448 iovss.n391 9.0005
R4962 iovss.n414 iovss.n391 9.0005
R4963 iovss.n449 iovss.n391 9.0005
R4964 iovss.n413 iovss.n391 9.0005
R4965 iovss.n451 iovss.n391 9.0005
R4966 iovss.n412 iovss.n391 9.0005
R4967 iovss.n3339 iovss.n391 9.0005
R4968 iovss.n3341 iovss.n391 9.0005
R4969 iovss.n3333 iovss.n391 9.0005
R4970 iovss.n3343 iovss.n386 9.0005
R4971 iovss.n429 iovss.n386 9.0005
R4972 iovss.n428 iovss.n386 9.0005
R4973 iovss.n431 iovss.n386 9.0005
R4974 iovss.n427 iovss.n386 9.0005
R4975 iovss.n432 iovss.n386 9.0005
R4976 iovss.n426 iovss.n386 9.0005
R4977 iovss.n434 iovss.n386 9.0005
R4978 iovss.n425 iovss.n386 9.0005
R4979 iovss.n435 iovss.n386 9.0005
R4980 iovss.n424 iovss.n386 9.0005
R4981 iovss.n437 iovss.n386 9.0005
R4982 iovss.n423 iovss.n386 9.0005
R4983 iovss.n386 iovss.n373 9.0005
R4984 iovss.n422 iovss.n386 9.0005
R4985 iovss.n439 iovss.n386 9.0005
R4986 iovss.n420 iovss.n386 9.0005
R4987 iovss.n440 iovss.n386 9.0005
R4988 iovss.n419 iovss.n386 9.0005
R4989 iovss.n442 iovss.n386 9.0005
R4990 iovss.n418 iovss.n386 9.0005
R4991 iovss.n443 iovss.n386 9.0005
R4992 iovss.n417 iovss.n386 9.0005
R4993 iovss.n445 iovss.n386 9.0005
R4994 iovss.n416 iovss.n386 9.0005
R4995 iovss.n446 iovss.n386 9.0005
R4996 iovss.n415 iovss.n386 9.0005
R4997 iovss.n448 iovss.n386 9.0005
R4998 iovss.n414 iovss.n386 9.0005
R4999 iovss.n449 iovss.n386 9.0005
R5000 iovss.n413 iovss.n386 9.0005
R5001 iovss.n451 iovss.n386 9.0005
R5002 iovss.n412 iovss.n386 9.0005
R5003 iovss.n3339 iovss.n386 9.0005
R5004 iovss.n3341 iovss.n386 9.0005
R5005 iovss.n3333 iovss.n386 9.0005
R5006 iovss.n3343 iovss.n393 9.0005
R5007 iovss.n429 iovss.n393 9.0005
R5008 iovss.n428 iovss.n393 9.0005
R5009 iovss.n431 iovss.n393 9.0005
R5010 iovss.n427 iovss.n393 9.0005
R5011 iovss.n432 iovss.n393 9.0005
R5012 iovss.n426 iovss.n393 9.0005
R5013 iovss.n434 iovss.n393 9.0005
R5014 iovss.n425 iovss.n393 9.0005
R5015 iovss.n435 iovss.n393 9.0005
R5016 iovss.n424 iovss.n393 9.0005
R5017 iovss.n437 iovss.n393 9.0005
R5018 iovss.n423 iovss.n393 9.0005
R5019 iovss.n393 iovss.n373 9.0005
R5020 iovss.n422 iovss.n393 9.0005
R5021 iovss.n439 iovss.n393 9.0005
R5022 iovss.n420 iovss.n393 9.0005
R5023 iovss.n440 iovss.n393 9.0005
R5024 iovss.n419 iovss.n393 9.0005
R5025 iovss.n442 iovss.n393 9.0005
R5026 iovss.n418 iovss.n393 9.0005
R5027 iovss.n443 iovss.n393 9.0005
R5028 iovss.n417 iovss.n393 9.0005
R5029 iovss.n445 iovss.n393 9.0005
R5030 iovss.n416 iovss.n393 9.0005
R5031 iovss.n446 iovss.n393 9.0005
R5032 iovss.n415 iovss.n393 9.0005
R5033 iovss.n448 iovss.n393 9.0005
R5034 iovss.n414 iovss.n393 9.0005
R5035 iovss.n449 iovss.n393 9.0005
R5036 iovss.n413 iovss.n393 9.0005
R5037 iovss.n451 iovss.n393 9.0005
R5038 iovss.n412 iovss.n393 9.0005
R5039 iovss.n3339 iovss.n393 9.0005
R5040 iovss.n3341 iovss.n393 9.0005
R5041 iovss.n3333 iovss.n393 9.0005
R5042 iovss.n3343 iovss.n385 9.0005
R5043 iovss.n429 iovss.n385 9.0005
R5044 iovss.n428 iovss.n385 9.0005
R5045 iovss.n431 iovss.n385 9.0005
R5046 iovss.n427 iovss.n385 9.0005
R5047 iovss.n432 iovss.n385 9.0005
R5048 iovss.n426 iovss.n385 9.0005
R5049 iovss.n434 iovss.n385 9.0005
R5050 iovss.n425 iovss.n385 9.0005
R5051 iovss.n435 iovss.n385 9.0005
R5052 iovss.n424 iovss.n385 9.0005
R5053 iovss.n437 iovss.n385 9.0005
R5054 iovss.n423 iovss.n385 9.0005
R5055 iovss.n385 iovss.n373 9.0005
R5056 iovss.n422 iovss.n385 9.0005
R5057 iovss.n439 iovss.n385 9.0005
R5058 iovss.n420 iovss.n385 9.0005
R5059 iovss.n440 iovss.n385 9.0005
R5060 iovss.n419 iovss.n385 9.0005
R5061 iovss.n442 iovss.n385 9.0005
R5062 iovss.n418 iovss.n385 9.0005
R5063 iovss.n443 iovss.n385 9.0005
R5064 iovss.n417 iovss.n385 9.0005
R5065 iovss.n445 iovss.n385 9.0005
R5066 iovss.n416 iovss.n385 9.0005
R5067 iovss.n446 iovss.n385 9.0005
R5068 iovss.n415 iovss.n385 9.0005
R5069 iovss.n448 iovss.n385 9.0005
R5070 iovss.n414 iovss.n385 9.0005
R5071 iovss.n449 iovss.n385 9.0005
R5072 iovss.n413 iovss.n385 9.0005
R5073 iovss.n451 iovss.n385 9.0005
R5074 iovss.n412 iovss.n385 9.0005
R5075 iovss.n3339 iovss.n385 9.0005
R5076 iovss.n3341 iovss.n385 9.0005
R5077 iovss.n3333 iovss.n385 9.0005
R5078 iovss.n3343 iovss.n395 9.0005
R5079 iovss.n429 iovss.n395 9.0005
R5080 iovss.n428 iovss.n395 9.0005
R5081 iovss.n431 iovss.n395 9.0005
R5082 iovss.n427 iovss.n395 9.0005
R5083 iovss.n432 iovss.n395 9.0005
R5084 iovss.n426 iovss.n395 9.0005
R5085 iovss.n434 iovss.n395 9.0005
R5086 iovss.n425 iovss.n395 9.0005
R5087 iovss.n435 iovss.n395 9.0005
R5088 iovss.n424 iovss.n395 9.0005
R5089 iovss.n437 iovss.n395 9.0005
R5090 iovss.n423 iovss.n395 9.0005
R5091 iovss.n395 iovss.n373 9.0005
R5092 iovss.n422 iovss.n395 9.0005
R5093 iovss.n439 iovss.n395 9.0005
R5094 iovss.n420 iovss.n395 9.0005
R5095 iovss.n440 iovss.n395 9.0005
R5096 iovss.n419 iovss.n395 9.0005
R5097 iovss.n442 iovss.n395 9.0005
R5098 iovss.n418 iovss.n395 9.0005
R5099 iovss.n443 iovss.n395 9.0005
R5100 iovss.n417 iovss.n395 9.0005
R5101 iovss.n445 iovss.n395 9.0005
R5102 iovss.n416 iovss.n395 9.0005
R5103 iovss.n446 iovss.n395 9.0005
R5104 iovss.n415 iovss.n395 9.0005
R5105 iovss.n448 iovss.n395 9.0005
R5106 iovss.n414 iovss.n395 9.0005
R5107 iovss.n449 iovss.n395 9.0005
R5108 iovss.n413 iovss.n395 9.0005
R5109 iovss.n451 iovss.n395 9.0005
R5110 iovss.n412 iovss.n395 9.0005
R5111 iovss.n3339 iovss.n395 9.0005
R5112 iovss.n3341 iovss.n395 9.0005
R5113 iovss.n3333 iovss.n395 9.0005
R5114 iovss.n3343 iovss.n384 9.0005
R5115 iovss.n429 iovss.n384 9.0005
R5116 iovss.n428 iovss.n384 9.0005
R5117 iovss.n431 iovss.n384 9.0005
R5118 iovss.n427 iovss.n384 9.0005
R5119 iovss.n432 iovss.n384 9.0005
R5120 iovss.n426 iovss.n384 9.0005
R5121 iovss.n434 iovss.n384 9.0005
R5122 iovss.n425 iovss.n384 9.0005
R5123 iovss.n435 iovss.n384 9.0005
R5124 iovss.n424 iovss.n384 9.0005
R5125 iovss.n437 iovss.n384 9.0005
R5126 iovss.n423 iovss.n384 9.0005
R5127 iovss.n384 iovss.n373 9.0005
R5128 iovss.n422 iovss.n384 9.0005
R5129 iovss.n439 iovss.n384 9.0005
R5130 iovss.n420 iovss.n384 9.0005
R5131 iovss.n440 iovss.n384 9.0005
R5132 iovss.n419 iovss.n384 9.0005
R5133 iovss.n442 iovss.n384 9.0005
R5134 iovss.n418 iovss.n384 9.0005
R5135 iovss.n443 iovss.n384 9.0005
R5136 iovss.n417 iovss.n384 9.0005
R5137 iovss.n445 iovss.n384 9.0005
R5138 iovss.n416 iovss.n384 9.0005
R5139 iovss.n446 iovss.n384 9.0005
R5140 iovss.n415 iovss.n384 9.0005
R5141 iovss.n448 iovss.n384 9.0005
R5142 iovss.n414 iovss.n384 9.0005
R5143 iovss.n449 iovss.n384 9.0005
R5144 iovss.n413 iovss.n384 9.0005
R5145 iovss.n451 iovss.n384 9.0005
R5146 iovss.n412 iovss.n384 9.0005
R5147 iovss.n3339 iovss.n384 9.0005
R5148 iovss.n3341 iovss.n384 9.0005
R5149 iovss.n3333 iovss.n384 9.0005
R5150 iovss.n3343 iovss.n397 9.0005
R5151 iovss.n429 iovss.n397 9.0005
R5152 iovss.n428 iovss.n397 9.0005
R5153 iovss.n431 iovss.n397 9.0005
R5154 iovss.n427 iovss.n397 9.0005
R5155 iovss.n432 iovss.n397 9.0005
R5156 iovss.n426 iovss.n397 9.0005
R5157 iovss.n434 iovss.n397 9.0005
R5158 iovss.n425 iovss.n397 9.0005
R5159 iovss.n435 iovss.n397 9.0005
R5160 iovss.n424 iovss.n397 9.0005
R5161 iovss.n437 iovss.n397 9.0005
R5162 iovss.n423 iovss.n397 9.0005
R5163 iovss.n397 iovss.n373 9.0005
R5164 iovss.n422 iovss.n397 9.0005
R5165 iovss.n439 iovss.n397 9.0005
R5166 iovss.n420 iovss.n397 9.0005
R5167 iovss.n440 iovss.n397 9.0005
R5168 iovss.n419 iovss.n397 9.0005
R5169 iovss.n442 iovss.n397 9.0005
R5170 iovss.n418 iovss.n397 9.0005
R5171 iovss.n443 iovss.n397 9.0005
R5172 iovss.n417 iovss.n397 9.0005
R5173 iovss.n445 iovss.n397 9.0005
R5174 iovss.n416 iovss.n397 9.0005
R5175 iovss.n446 iovss.n397 9.0005
R5176 iovss.n415 iovss.n397 9.0005
R5177 iovss.n448 iovss.n397 9.0005
R5178 iovss.n414 iovss.n397 9.0005
R5179 iovss.n449 iovss.n397 9.0005
R5180 iovss.n413 iovss.n397 9.0005
R5181 iovss.n451 iovss.n397 9.0005
R5182 iovss.n412 iovss.n397 9.0005
R5183 iovss.n3339 iovss.n397 9.0005
R5184 iovss.n3341 iovss.n397 9.0005
R5185 iovss.n3333 iovss.n397 9.0005
R5186 iovss.n3343 iovss.n383 9.0005
R5187 iovss.n429 iovss.n383 9.0005
R5188 iovss.n428 iovss.n383 9.0005
R5189 iovss.n431 iovss.n383 9.0005
R5190 iovss.n427 iovss.n383 9.0005
R5191 iovss.n432 iovss.n383 9.0005
R5192 iovss.n426 iovss.n383 9.0005
R5193 iovss.n434 iovss.n383 9.0005
R5194 iovss.n425 iovss.n383 9.0005
R5195 iovss.n435 iovss.n383 9.0005
R5196 iovss.n424 iovss.n383 9.0005
R5197 iovss.n437 iovss.n383 9.0005
R5198 iovss.n423 iovss.n383 9.0005
R5199 iovss.n383 iovss.n373 9.0005
R5200 iovss.n422 iovss.n383 9.0005
R5201 iovss.n439 iovss.n383 9.0005
R5202 iovss.n420 iovss.n383 9.0005
R5203 iovss.n440 iovss.n383 9.0005
R5204 iovss.n419 iovss.n383 9.0005
R5205 iovss.n442 iovss.n383 9.0005
R5206 iovss.n418 iovss.n383 9.0005
R5207 iovss.n443 iovss.n383 9.0005
R5208 iovss.n417 iovss.n383 9.0005
R5209 iovss.n445 iovss.n383 9.0005
R5210 iovss.n416 iovss.n383 9.0005
R5211 iovss.n446 iovss.n383 9.0005
R5212 iovss.n415 iovss.n383 9.0005
R5213 iovss.n448 iovss.n383 9.0005
R5214 iovss.n414 iovss.n383 9.0005
R5215 iovss.n449 iovss.n383 9.0005
R5216 iovss.n413 iovss.n383 9.0005
R5217 iovss.n451 iovss.n383 9.0005
R5218 iovss.n412 iovss.n383 9.0005
R5219 iovss.n3339 iovss.n383 9.0005
R5220 iovss.n3341 iovss.n383 9.0005
R5221 iovss.n3333 iovss.n383 9.0005
R5222 iovss.n3343 iovss.n399 9.0005
R5223 iovss.n429 iovss.n399 9.0005
R5224 iovss.n428 iovss.n399 9.0005
R5225 iovss.n431 iovss.n399 9.0005
R5226 iovss.n427 iovss.n399 9.0005
R5227 iovss.n432 iovss.n399 9.0005
R5228 iovss.n426 iovss.n399 9.0005
R5229 iovss.n434 iovss.n399 9.0005
R5230 iovss.n425 iovss.n399 9.0005
R5231 iovss.n435 iovss.n399 9.0005
R5232 iovss.n424 iovss.n399 9.0005
R5233 iovss.n437 iovss.n399 9.0005
R5234 iovss.n423 iovss.n399 9.0005
R5235 iovss.n399 iovss.n373 9.0005
R5236 iovss.n422 iovss.n399 9.0005
R5237 iovss.n439 iovss.n399 9.0005
R5238 iovss.n420 iovss.n399 9.0005
R5239 iovss.n440 iovss.n399 9.0005
R5240 iovss.n419 iovss.n399 9.0005
R5241 iovss.n442 iovss.n399 9.0005
R5242 iovss.n418 iovss.n399 9.0005
R5243 iovss.n443 iovss.n399 9.0005
R5244 iovss.n417 iovss.n399 9.0005
R5245 iovss.n445 iovss.n399 9.0005
R5246 iovss.n416 iovss.n399 9.0005
R5247 iovss.n446 iovss.n399 9.0005
R5248 iovss.n415 iovss.n399 9.0005
R5249 iovss.n448 iovss.n399 9.0005
R5250 iovss.n414 iovss.n399 9.0005
R5251 iovss.n449 iovss.n399 9.0005
R5252 iovss.n413 iovss.n399 9.0005
R5253 iovss.n451 iovss.n399 9.0005
R5254 iovss.n412 iovss.n399 9.0005
R5255 iovss.n3339 iovss.n399 9.0005
R5256 iovss.n3341 iovss.n399 9.0005
R5257 iovss.n3333 iovss.n399 9.0005
R5258 iovss.n3343 iovss.n382 9.0005
R5259 iovss.n429 iovss.n382 9.0005
R5260 iovss.n428 iovss.n382 9.0005
R5261 iovss.n431 iovss.n382 9.0005
R5262 iovss.n427 iovss.n382 9.0005
R5263 iovss.n432 iovss.n382 9.0005
R5264 iovss.n426 iovss.n382 9.0005
R5265 iovss.n434 iovss.n382 9.0005
R5266 iovss.n425 iovss.n382 9.0005
R5267 iovss.n435 iovss.n382 9.0005
R5268 iovss.n424 iovss.n382 9.0005
R5269 iovss.n437 iovss.n382 9.0005
R5270 iovss.n423 iovss.n382 9.0005
R5271 iovss.n382 iovss.n373 9.0005
R5272 iovss.n422 iovss.n382 9.0005
R5273 iovss.n439 iovss.n382 9.0005
R5274 iovss.n420 iovss.n382 9.0005
R5275 iovss.n440 iovss.n382 9.0005
R5276 iovss.n419 iovss.n382 9.0005
R5277 iovss.n442 iovss.n382 9.0005
R5278 iovss.n418 iovss.n382 9.0005
R5279 iovss.n443 iovss.n382 9.0005
R5280 iovss.n417 iovss.n382 9.0005
R5281 iovss.n445 iovss.n382 9.0005
R5282 iovss.n416 iovss.n382 9.0005
R5283 iovss.n446 iovss.n382 9.0005
R5284 iovss.n415 iovss.n382 9.0005
R5285 iovss.n448 iovss.n382 9.0005
R5286 iovss.n414 iovss.n382 9.0005
R5287 iovss.n449 iovss.n382 9.0005
R5288 iovss.n413 iovss.n382 9.0005
R5289 iovss.n451 iovss.n382 9.0005
R5290 iovss.n412 iovss.n382 9.0005
R5291 iovss.n3339 iovss.n382 9.0005
R5292 iovss.n3341 iovss.n382 9.0005
R5293 iovss.n3333 iovss.n382 9.0005
R5294 iovss.n3343 iovss.n401 9.0005
R5295 iovss.n429 iovss.n401 9.0005
R5296 iovss.n428 iovss.n401 9.0005
R5297 iovss.n431 iovss.n401 9.0005
R5298 iovss.n427 iovss.n401 9.0005
R5299 iovss.n432 iovss.n401 9.0005
R5300 iovss.n426 iovss.n401 9.0005
R5301 iovss.n434 iovss.n401 9.0005
R5302 iovss.n425 iovss.n401 9.0005
R5303 iovss.n435 iovss.n401 9.0005
R5304 iovss.n424 iovss.n401 9.0005
R5305 iovss.n437 iovss.n401 9.0005
R5306 iovss.n423 iovss.n401 9.0005
R5307 iovss.n401 iovss.n373 9.0005
R5308 iovss.n422 iovss.n401 9.0005
R5309 iovss.n439 iovss.n401 9.0005
R5310 iovss.n420 iovss.n401 9.0005
R5311 iovss.n440 iovss.n401 9.0005
R5312 iovss.n419 iovss.n401 9.0005
R5313 iovss.n442 iovss.n401 9.0005
R5314 iovss.n418 iovss.n401 9.0005
R5315 iovss.n443 iovss.n401 9.0005
R5316 iovss.n417 iovss.n401 9.0005
R5317 iovss.n445 iovss.n401 9.0005
R5318 iovss.n416 iovss.n401 9.0005
R5319 iovss.n446 iovss.n401 9.0005
R5320 iovss.n415 iovss.n401 9.0005
R5321 iovss.n448 iovss.n401 9.0005
R5322 iovss.n414 iovss.n401 9.0005
R5323 iovss.n449 iovss.n401 9.0005
R5324 iovss.n413 iovss.n401 9.0005
R5325 iovss.n451 iovss.n401 9.0005
R5326 iovss.n412 iovss.n401 9.0005
R5327 iovss.n3339 iovss.n401 9.0005
R5328 iovss.n3341 iovss.n401 9.0005
R5329 iovss.n3333 iovss.n401 9.0005
R5330 iovss.n3343 iovss.n381 9.0005
R5331 iovss.n429 iovss.n381 9.0005
R5332 iovss.n428 iovss.n381 9.0005
R5333 iovss.n431 iovss.n381 9.0005
R5334 iovss.n427 iovss.n381 9.0005
R5335 iovss.n432 iovss.n381 9.0005
R5336 iovss.n426 iovss.n381 9.0005
R5337 iovss.n434 iovss.n381 9.0005
R5338 iovss.n425 iovss.n381 9.0005
R5339 iovss.n435 iovss.n381 9.0005
R5340 iovss.n424 iovss.n381 9.0005
R5341 iovss.n437 iovss.n381 9.0005
R5342 iovss.n423 iovss.n381 9.0005
R5343 iovss.n381 iovss.n373 9.0005
R5344 iovss.n422 iovss.n381 9.0005
R5345 iovss.n439 iovss.n381 9.0005
R5346 iovss.n420 iovss.n381 9.0005
R5347 iovss.n440 iovss.n381 9.0005
R5348 iovss.n419 iovss.n381 9.0005
R5349 iovss.n442 iovss.n381 9.0005
R5350 iovss.n418 iovss.n381 9.0005
R5351 iovss.n443 iovss.n381 9.0005
R5352 iovss.n417 iovss.n381 9.0005
R5353 iovss.n445 iovss.n381 9.0005
R5354 iovss.n416 iovss.n381 9.0005
R5355 iovss.n446 iovss.n381 9.0005
R5356 iovss.n415 iovss.n381 9.0005
R5357 iovss.n448 iovss.n381 9.0005
R5358 iovss.n414 iovss.n381 9.0005
R5359 iovss.n449 iovss.n381 9.0005
R5360 iovss.n413 iovss.n381 9.0005
R5361 iovss.n451 iovss.n381 9.0005
R5362 iovss.n412 iovss.n381 9.0005
R5363 iovss.n3339 iovss.n381 9.0005
R5364 iovss.n3341 iovss.n381 9.0005
R5365 iovss.n3333 iovss.n381 9.0005
R5366 iovss.n3343 iovss.n3342 9.0005
R5367 iovss.n3342 iovss.n429 9.0005
R5368 iovss.n3342 iovss.n428 9.0005
R5369 iovss.n3342 iovss.n431 9.0005
R5370 iovss.n3342 iovss.n427 9.0005
R5371 iovss.n3342 iovss.n432 9.0005
R5372 iovss.n3342 iovss.n426 9.0005
R5373 iovss.n3342 iovss.n434 9.0005
R5374 iovss.n3342 iovss.n425 9.0005
R5375 iovss.n3342 iovss.n435 9.0005
R5376 iovss.n3342 iovss.n424 9.0005
R5377 iovss.n3342 iovss.n437 9.0005
R5378 iovss.n3342 iovss.n423 9.0005
R5379 iovss.n3342 iovss.n373 9.0005
R5380 iovss.n3342 iovss.n422 9.0005
R5381 iovss.n3342 iovss.n439 9.0005
R5382 iovss.n3342 iovss.n420 9.0005
R5383 iovss.n3342 iovss.n440 9.0005
R5384 iovss.n3342 iovss.n419 9.0005
R5385 iovss.n3342 iovss.n442 9.0005
R5386 iovss.n3342 iovss.n418 9.0005
R5387 iovss.n3342 iovss.n443 9.0005
R5388 iovss.n3342 iovss.n417 9.0005
R5389 iovss.n3342 iovss.n445 9.0005
R5390 iovss.n3342 iovss.n416 9.0005
R5391 iovss.n3342 iovss.n446 9.0005
R5392 iovss.n3342 iovss.n415 9.0005
R5393 iovss.n3342 iovss.n448 9.0005
R5394 iovss.n3342 iovss.n414 9.0005
R5395 iovss.n3342 iovss.n449 9.0005
R5396 iovss.n3342 iovss.n413 9.0005
R5397 iovss.n3342 iovss.n451 9.0005
R5398 iovss.n3342 iovss.n412 9.0005
R5399 iovss.n3342 iovss.n3339 9.0005
R5400 iovss.n3342 iovss.n3341 9.0005
R5401 iovss.n3478 iovss.n8 9.0005
R5402 iovss.n19 iovss.n8 9.0005
R5403 iovss.n52 iovss.n8 9.0005
R5404 iovss.n17 iovss.n8 9.0005
R5405 iovss.n55 iovss.n8 9.0005
R5406 iovss.n3480 iovss.n8 9.0005
R5407 iovss.n3478 iovss.n7 9.0005
R5408 iovss.n20 iovss.n7 9.0005
R5409 iovss.n51 iovss.n7 9.0005
R5410 iovss.n19 iovss.n7 9.0005
R5411 iovss.n52 iovss.n7 9.0005
R5412 iovss.n18 iovss.n7 9.0005
R5413 iovss.n54 iovss.n7 9.0005
R5414 iovss.n17 iovss.n7 9.0005
R5415 iovss.n55 iovss.n7 9.0005
R5416 iovss.n16 iovss.n7 9.0005
R5417 iovss.n57 iovss.n7 9.0005
R5418 iovss.n3480 iovss.n7 9.0005
R5419 iovss.n3478 iovss.n9 9.0005
R5420 iovss.n20 iovss.n9 9.0005
R5421 iovss.n51 iovss.n9 9.0005
R5422 iovss.n19 iovss.n9 9.0005
R5423 iovss.n52 iovss.n9 9.0005
R5424 iovss.n18 iovss.n9 9.0005
R5425 iovss.n54 iovss.n9 9.0005
R5426 iovss.n17 iovss.n9 9.0005
R5427 iovss.n55 iovss.n9 9.0005
R5428 iovss.n16 iovss.n9 9.0005
R5429 iovss.n57 iovss.n9 9.0005
R5430 iovss.n3480 iovss.n9 9.0005
R5431 iovss.n3478 iovss.n6 9.0005
R5432 iovss.n20 iovss.n6 9.0005
R5433 iovss.n51 iovss.n6 9.0005
R5434 iovss.n19 iovss.n6 9.0005
R5435 iovss.n52 iovss.n6 9.0005
R5436 iovss.n18 iovss.n6 9.0005
R5437 iovss.n54 iovss.n6 9.0005
R5438 iovss.n17 iovss.n6 9.0005
R5439 iovss.n55 iovss.n6 9.0005
R5440 iovss.n16 iovss.n6 9.0005
R5441 iovss.n57 iovss.n6 9.0005
R5442 iovss.n3480 iovss.n6 9.0005
R5443 iovss.n3478 iovss.n10 9.0005
R5444 iovss.n20 iovss.n10 9.0005
R5445 iovss.n51 iovss.n10 9.0005
R5446 iovss.n19 iovss.n10 9.0005
R5447 iovss.n52 iovss.n10 9.0005
R5448 iovss.n18 iovss.n10 9.0005
R5449 iovss.n54 iovss.n10 9.0005
R5450 iovss.n17 iovss.n10 9.0005
R5451 iovss.n55 iovss.n10 9.0005
R5452 iovss.n16 iovss.n10 9.0005
R5453 iovss.n57 iovss.n10 9.0005
R5454 iovss.n3480 iovss.n10 9.0005
R5455 iovss.n3478 iovss.n5 9.0005
R5456 iovss.n20 iovss.n5 9.0005
R5457 iovss.n51 iovss.n5 9.0005
R5458 iovss.n19 iovss.n5 9.0005
R5459 iovss.n52 iovss.n5 9.0005
R5460 iovss.n18 iovss.n5 9.0005
R5461 iovss.n54 iovss.n5 9.0005
R5462 iovss.n17 iovss.n5 9.0005
R5463 iovss.n55 iovss.n5 9.0005
R5464 iovss.n16 iovss.n5 9.0005
R5465 iovss.n57 iovss.n5 9.0005
R5466 iovss.n3480 iovss.n5 9.0005
R5467 iovss.n3478 iovss.n11 9.0005
R5468 iovss.n20 iovss.n11 9.0005
R5469 iovss.n51 iovss.n11 9.0005
R5470 iovss.n19 iovss.n11 9.0005
R5471 iovss.n52 iovss.n11 9.0005
R5472 iovss.n18 iovss.n11 9.0005
R5473 iovss.n54 iovss.n11 9.0005
R5474 iovss.n17 iovss.n11 9.0005
R5475 iovss.n55 iovss.n11 9.0005
R5476 iovss.n16 iovss.n11 9.0005
R5477 iovss.n57 iovss.n11 9.0005
R5478 iovss.n3480 iovss.n11 9.0005
R5479 iovss.n3478 iovss.n4 9.0005
R5480 iovss.n20 iovss.n4 9.0005
R5481 iovss.n51 iovss.n4 9.0005
R5482 iovss.n19 iovss.n4 9.0005
R5483 iovss.n52 iovss.n4 9.0005
R5484 iovss.n18 iovss.n4 9.0005
R5485 iovss.n54 iovss.n4 9.0005
R5486 iovss.n17 iovss.n4 9.0005
R5487 iovss.n55 iovss.n4 9.0005
R5488 iovss.n16 iovss.n4 9.0005
R5489 iovss.n57 iovss.n4 9.0005
R5490 iovss.n3480 iovss.n4 9.0005
R5491 iovss.n3478 iovss.n12 9.0005
R5492 iovss.n20 iovss.n12 9.0005
R5493 iovss.n51 iovss.n12 9.0005
R5494 iovss.n19 iovss.n12 9.0005
R5495 iovss.n52 iovss.n12 9.0005
R5496 iovss.n18 iovss.n12 9.0005
R5497 iovss.n54 iovss.n12 9.0005
R5498 iovss.n17 iovss.n12 9.0005
R5499 iovss.n55 iovss.n12 9.0005
R5500 iovss.n16 iovss.n12 9.0005
R5501 iovss.n57 iovss.n12 9.0005
R5502 iovss.n3480 iovss.n12 9.0005
R5503 iovss.n3478 iovss.n3 9.0005
R5504 iovss.n20 iovss.n3 9.0005
R5505 iovss.n51 iovss.n3 9.0005
R5506 iovss.n19 iovss.n3 9.0005
R5507 iovss.n52 iovss.n3 9.0005
R5508 iovss.n18 iovss.n3 9.0005
R5509 iovss.n54 iovss.n3 9.0005
R5510 iovss.n17 iovss.n3 9.0005
R5511 iovss.n55 iovss.n3 9.0005
R5512 iovss.n16 iovss.n3 9.0005
R5513 iovss.n57 iovss.n3 9.0005
R5514 iovss.n3480 iovss.n3 9.0005
R5515 iovss.n3478 iovss.n13 9.0005
R5516 iovss.n20 iovss.n13 9.0005
R5517 iovss.n51 iovss.n13 9.0005
R5518 iovss.n19 iovss.n13 9.0005
R5519 iovss.n52 iovss.n13 9.0005
R5520 iovss.n18 iovss.n13 9.0005
R5521 iovss.n54 iovss.n13 9.0005
R5522 iovss.n17 iovss.n13 9.0005
R5523 iovss.n55 iovss.n13 9.0005
R5524 iovss.n16 iovss.n13 9.0005
R5525 iovss.n57 iovss.n13 9.0005
R5526 iovss.n3480 iovss.n13 9.0005
R5527 iovss.n3478 iovss.n2 9.0005
R5528 iovss.n20 iovss.n2 9.0005
R5529 iovss.n51 iovss.n2 9.0005
R5530 iovss.n19 iovss.n2 9.0005
R5531 iovss.n52 iovss.n2 9.0005
R5532 iovss.n18 iovss.n2 9.0005
R5533 iovss.n54 iovss.n2 9.0005
R5534 iovss.n17 iovss.n2 9.0005
R5535 iovss.n55 iovss.n2 9.0005
R5536 iovss.n16 iovss.n2 9.0005
R5537 iovss.n57 iovss.n2 9.0005
R5538 iovss.n3480 iovss.n2 9.0005
R5539 iovss.n3478 iovss.n14 9.0005
R5540 iovss.n20 iovss.n14 9.0005
R5541 iovss.n51 iovss.n14 9.0005
R5542 iovss.n19 iovss.n14 9.0005
R5543 iovss.n52 iovss.n14 9.0005
R5544 iovss.n18 iovss.n14 9.0005
R5545 iovss.n54 iovss.n14 9.0005
R5546 iovss.n17 iovss.n14 9.0005
R5547 iovss.n55 iovss.n14 9.0005
R5548 iovss.n16 iovss.n14 9.0005
R5549 iovss.n57 iovss.n14 9.0005
R5550 iovss.n3480 iovss.n14 9.0005
R5551 iovss.n3478 iovss.n1 9.0005
R5552 iovss.n20 iovss.n1 9.0005
R5553 iovss.n51 iovss.n1 9.0005
R5554 iovss.n19 iovss.n1 9.0005
R5555 iovss.n52 iovss.n1 9.0005
R5556 iovss.n18 iovss.n1 9.0005
R5557 iovss.n54 iovss.n1 9.0005
R5558 iovss.n17 iovss.n1 9.0005
R5559 iovss.n55 iovss.n1 9.0005
R5560 iovss.n16 iovss.n1 9.0005
R5561 iovss.n57 iovss.n1 9.0005
R5562 iovss.n3480 iovss.n1 9.0005
R5563 iovss.n3479 iovss.n20 9.0005
R5564 iovss.n3479 iovss.n51 9.0005
R5565 iovss.n3479 iovss.n19 9.0005
R5566 iovss.n3479 iovss.n52 9.0005
R5567 iovss.n3479 iovss.n18 9.0005
R5568 iovss.n3479 iovss.n54 9.0005
R5569 iovss.n3479 iovss.n17 9.0005
R5570 iovss.n3479 iovss.n55 9.0005
R5571 iovss.n3479 iovss.n16 9.0005
R5572 iovss.n3479 iovss.n57 9.0005
R5573 iovss.n3480 iovss.n3479 9.0005
R5574 iovss.n3479 iovss.n3478 9.0005
R5575 iovss.n3432 iovss.n171 9.0005
R5576 iovss.n3432 iovss.n122 9.0005
R5577 iovss.n3432 iovss.n117 9.0005
R5578 iovss.n3432 iovss.n126 9.0005
R5579 iovss.n3432 iovss.n115 9.0005
R5580 iovss.n3434 iovss.n3432 9.0005
R5581 iovss.n3432 iovss.n68 9.0005
R5582 iovss.n111 iovss.n87 9.0005
R5583 iovss.n135 iovss.n87 9.0005
R5584 iovss.n109 iovss.n87 9.0005
R5585 iovss.n138 iovss.n87 9.0005
R5586 iovss.n107 iovss.n87 9.0005
R5587 iovss.n141 iovss.n87 9.0005
R5588 iovss.n105 iovss.n87 9.0005
R5589 iovss.n145 iovss.n87 9.0005
R5590 iovss.n87 iovss.n78 9.0005
R5591 iovss.n3436 iovss.n87 9.0005
R5592 iovss.n3434 iovss.n87 9.0005
R5593 iovss.n87 iovss.n68 9.0005
R5594 iovss.n120 iovss.n85 9.0005
R5595 iovss.n118 iovss.n85 9.0005
R5596 iovss.n122 iovss.n85 9.0005
R5597 iovss.n117 iovss.n85 9.0005
R5598 iovss.n124 iovss.n85 9.0005
R5599 iovss.n116 iovss.n85 9.0005
R5600 iovss.n126 iovss.n85 9.0005
R5601 iovss.n115 iovss.n85 9.0005
R5602 iovss.n128 iovss.n85 9.0005
R5603 iovss.n114 iovss.n85 9.0005
R5604 iovss.n130 iovss.n85 9.0005
R5605 iovss.n113 iovss.n85 9.0005
R5606 iovss.n132 iovss.n85 9.0005
R5607 iovss.n112 iovss.n85 9.0005
R5608 iovss.n134 iovss.n85 9.0005
R5609 iovss.n111 iovss.n85 9.0005
R5610 iovss.n135 iovss.n85 9.0005
R5611 iovss.n110 iovss.n85 9.0005
R5612 iovss.n137 iovss.n85 9.0005
R5613 iovss.n109 iovss.n85 9.0005
R5614 iovss.n138 iovss.n85 9.0005
R5615 iovss.n108 iovss.n85 9.0005
R5616 iovss.n140 iovss.n85 9.0005
R5617 iovss.n107 iovss.n85 9.0005
R5618 iovss.n141 iovss.n85 9.0005
R5619 iovss.n106 iovss.n85 9.0005
R5620 iovss.n143 iovss.n85 9.0005
R5621 iovss.n105 iovss.n85 9.0005
R5622 iovss.n145 iovss.n85 9.0005
R5623 iovss.n104 iovss.n85 9.0005
R5624 iovss.n147 iovss.n85 9.0005
R5625 iovss.n85 iovss.n78 9.0005
R5626 iovss.n3436 iovss.n85 9.0005
R5627 iovss.n85 iovss.n68 9.0005
R5628 iovss.n120 iovss.n88 9.0005
R5629 iovss.n118 iovss.n88 9.0005
R5630 iovss.n122 iovss.n88 9.0005
R5631 iovss.n117 iovss.n88 9.0005
R5632 iovss.n124 iovss.n88 9.0005
R5633 iovss.n116 iovss.n88 9.0005
R5634 iovss.n126 iovss.n88 9.0005
R5635 iovss.n115 iovss.n88 9.0005
R5636 iovss.n128 iovss.n88 9.0005
R5637 iovss.n114 iovss.n88 9.0005
R5638 iovss.n130 iovss.n88 9.0005
R5639 iovss.n113 iovss.n88 9.0005
R5640 iovss.n132 iovss.n88 9.0005
R5641 iovss.n112 iovss.n88 9.0005
R5642 iovss.n134 iovss.n88 9.0005
R5643 iovss.n111 iovss.n88 9.0005
R5644 iovss.n135 iovss.n88 9.0005
R5645 iovss.n110 iovss.n88 9.0005
R5646 iovss.n137 iovss.n88 9.0005
R5647 iovss.n109 iovss.n88 9.0005
R5648 iovss.n138 iovss.n88 9.0005
R5649 iovss.n108 iovss.n88 9.0005
R5650 iovss.n140 iovss.n88 9.0005
R5651 iovss.n107 iovss.n88 9.0005
R5652 iovss.n141 iovss.n88 9.0005
R5653 iovss.n106 iovss.n88 9.0005
R5654 iovss.n143 iovss.n88 9.0005
R5655 iovss.n105 iovss.n88 9.0005
R5656 iovss.n145 iovss.n88 9.0005
R5657 iovss.n104 iovss.n88 9.0005
R5658 iovss.n147 iovss.n88 9.0005
R5659 iovss.n88 iovss.n78 9.0005
R5660 iovss.n3436 iovss.n88 9.0005
R5661 iovss.n88 iovss.n68 9.0005
R5662 iovss.n120 iovss.n84 9.0005
R5663 iovss.n118 iovss.n84 9.0005
R5664 iovss.n122 iovss.n84 9.0005
R5665 iovss.n117 iovss.n84 9.0005
R5666 iovss.n124 iovss.n84 9.0005
R5667 iovss.n116 iovss.n84 9.0005
R5668 iovss.n126 iovss.n84 9.0005
R5669 iovss.n115 iovss.n84 9.0005
R5670 iovss.n128 iovss.n84 9.0005
R5671 iovss.n114 iovss.n84 9.0005
R5672 iovss.n130 iovss.n84 9.0005
R5673 iovss.n113 iovss.n84 9.0005
R5674 iovss.n132 iovss.n84 9.0005
R5675 iovss.n112 iovss.n84 9.0005
R5676 iovss.n134 iovss.n84 9.0005
R5677 iovss.n111 iovss.n84 9.0005
R5678 iovss.n135 iovss.n84 9.0005
R5679 iovss.n110 iovss.n84 9.0005
R5680 iovss.n137 iovss.n84 9.0005
R5681 iovss.n109 iovss.n84 9.0005
R5682 iovss.n138 iovss.n84 9.0005
R5683 iovss.n108 iovss.n84 9.0005
R5684 iovss.n140 iovss.n84 9.0005
R5685 iovss.n107 iovss.n84 9.0005
R5686 iovss.n141 iovss.n84 9.0005
R5687 iovss.n106 iovss.n84 9.0005
R5688 iovss.n143 iovss.n84 9.0005
R5689 iovss.n105 iovss.n84 9.0005
R5690 iovss.n145 iovss.n84 9.0005
R5691 iovss.n104 iovss.n84 9.0005
R5692 iovss.n147 iovss.n84 9.0005
R5693 iovss.n84 iovss.n78 9.0005
R5694 iovss.n3436 iovss.n84 9.0005
R5695 iovss.n103 iovss.n84 9.0005
R5696 iovss.n3434 iovss.n84 9.0005
R5697 iovss.n84 iovss.n68 9.0005
R5698 iovss.n120 iovss.n89 9.0005
R5699 iovss.n118 iovss.n89 9.0005
R5700 iovss.n122 iovss.n89 9.0005
R5701 iovss.n117 iovss.n89 9.0005
R5702 iovss.n124 iovss.n89 9.0005
R5703 iovss.n116 iovss.n89 9.0005
R5704 iovss.n126 iovss.n89 9.0005
R5705 iovss.n115 iovss.n89 9.0005
R5706 iovss.n128 iovss.n89 9.0005
R5707 iovss.n114 iovss.n89 9.0005
R5708 iovss.n130 iovss.n89 9.0005
R5709 iovss.n113 iovss.n89 9.0005
R5710 iovss.n132 iovss.n89 9.0005
R5711 iovss.n112 iovss.n89 9.0005
R5712 iovss.n134 iovss.n89 9.0005
R5713 iovss.n111 iovss.n89 9.0005
R5714 iovss.n135 iovss.n89 9.0005
R5715 iovss.n110 iovss.n89 9.0005
R5716 iovss.n137 iovss.n89 9.0005
R5717 iovss.n109 iovss.n89 9.0005
R5718 iovss.n138 iovss.n89 9.0005
R5719 iovss.n108 iovss.n89 9.0005
R5720 iovss.n140 iovss.n89 9.0005
R5721 iovss.n107 iovss.n89 9.0005
R5722 iovss.n141 iovss.n89 9.0005
R5723 iovss.n106 iovss.n89 9.0005
R5724 iovss.n143 iovss.n89 9.0005
R5725 iovss.n105 iovss.n89 9.0005
R5726 iovss.n145 iovss.n89 9.0005
R5727 iovss.n104 iovss.n89 9.0005
R5728 iovss.n147 iovss.n89 9.0005
R5729 iovss.n89 iovss.n78 9.0005
R5730 iovss.n3436 iovss.n89 9.0005
R5731 iovss.n103 iovss.n89 9.0005
R5732 iovss.n3434 iovss.n89 9.0005
R5733 iovss.n89 iovss.n68 9.0005
R5734 iovss.n120 iovss.n83 9.0005
R5735 iovss.n118 iovss.n83 9.0005
R5736 iovss.n122 iovss.n83 9.0005
R5737 iovss.n117 iovss.n83 9.0005
R5738 iovss.n124 iovss.n83 9.0005
R5739 iovss.n116 iovss.n83 9.0005
R5740 iovss.n126 iovss.n83 9.0005
R5741 iovss.n115 iovss.n83 9.0005
R5742 iovss.n128 iovss.n83 9.0005
R5743 iovss.n114 iovss.n83 9.0005
R5744 iovss.n130 iovss.n83 9.0005
R5745 iovss.n113 iovss.n83 9.0005
R5746 iovss.n132 iovss.n83 9.0005
R5747 iovss.n112 iovss.n83 9.0005
R5748 iovss.n134 iovss.n83 9.0005
R5749 iovss.n111 iovss.n83 9.0005
R5750 iovss.n135 iovss.n83 9.0005
R5751 iovss.n110 iovss.n83 9.0005
R5752 iovss.n137 iovss.n83 9.0005
R5753 iovss.n109 iovss.n83 9.0005
R5754 iovss.n138 iovss.n83 9.0005
R5755 iovss.n108 iovss.n83 9.0005
R5756 iovss.n140 iovss.n83 9.0005
R5757 iovss.n107 iovss.n83 9.0005
R5758 iovss.n141 iovss.n83 9.0005
R5759 iovss.n106 iovss.n83 9.0005
R5760 iovss.n143 iovss.n83 9.0005
R5761 iovss.n105 iovss.n83 9.0005
R5762 iovss.n145 iovss.n83 9.0005
R5763 iovss.n104 iovss.n83 9.0005
R5764 iovss.n147 iovss.n83 9.0005
R5765 iovss.n83 iovss.n78 9.0005
R5766 iovss.n3436 iovss.n83 9.0005
R5767 iovss.n103 iovss.n83 9.0005
R5768 iovss.n3434 iovss.n83 9.0005
R5769 iovss.n83 iovss.n68 9.0005
R5770 iovss.n120 iovss.n90 9.0005
R5771 iovss.n118 iovss.n90 9.0005
R5772 iovss.n122 iovss.n90 9.0005
R5773 iovss.n117 iovss.n90 9.0005
R5774 iovss.n124 iovss.n90 9.0005
R5775 iovss.n116 iovss.n90 9.0005
R5776 iovss.n126 iovss.n90 9.0005
R5777 iovss.n115 iovss.n90 9.0005
R5778 iovss.n128 iovss.n90 9.0005
R5779 iovss.n114 iovss.n90 9.0005
R5780 iovss.n130 iovss.n90 9.0005
R5781 iovss.n113 iovss.n90 9.0005
R5782 iovss.n132 iovss.n90 9.0005
R5783 iovss.n112 iovss.n90 9.0005
R5784 iovss.n134 iovss.n90 9.0005
R5785 iovss.n111 iovss.n90 9.0005
R5786 iovss.n135 iovss.n90 9.0005
R5787 iovss.n110 iovss.n90 9.0005
R5788 iovss.n137 iovss.n90 9.0005
R5789 iovss.n109 iovss.n90 9.0005
R5790 iovss.n138 iovss.n90 9.0005
R5791 iovss.n108 iovss.n90 9.0005
R5792 iovss.n140 iovss.n90 9.0005
R5793 iovss.n107 iovss.n90 9.0005
R5794 iovss.n141 iovss.n90 9.0005
R5795 iovss.n106 iovss.n90 9.0005
R5796 iovss.n143 iovss.n90 9.0005
R5797 iovss.n105 iovss.n90 9.0005
R5798 iovss.n145 iovss.n90 9.0005
R5799 iovss.n104 iovss.n90 9.0005
R5800 iovss.n147 iovss.n90 9.0005
R5801 iovss.n90 iovss.n78 9.0005
R5802 iovss.n3436 iovss.n90 9.0005
R5803 iovss.n103 iovss.n90 9.0005
R5804 iovss.n3434 iovss.n90 9.0005
R5805 iovss.n90 iovss.n68 9.0005
R5806 iovss.n120 iovss.n82 9.0005
R5807 iovss.n118 iovss.n82 9.0005
R5808 iovss.n122 iovss.n82 9.0005
R5809 iovss.n117 iovss.n82 9.0005
R5810 iovss.n124 iovss.n82 9.0005
R5811 iovss.n116 iovss.n82 9.0005
R5812 iovss.n126 iovss.n82 9.0005
R5813 iovss.n115 iovss.n82 9.0005
R5814 iovss.n128 iovss.n82 9.0005
R5815 iovss.n114 iovss.n82 9.0005
R5816 iovss.n130 iovss.n82 9.0005
R5817 iovss.n113 iovss.n82 9.0005
R5818 iovss.n132 iovss.n82 9.0005
R5819 iovss.n112 iovss.n82 9.0005
R5820 iovss.n134 iovss.n82 9.0005
R5821 iovss.n111 iovss.n82 9.0005
R5822 iovss.n135 iovss.n82 9.0005
R5823 iovss.n110 iovss.n82 9.0005
R5824 iovss.n137 iovss.n82 9.0005
R5825 iovss.n109 iovss.n82 9.0005
R5826 iovss.n138 iovss.n82 9.0005
R5827 iovss.n108 iovss.n82 9.0005
R5828 iovss.n140 iovss.n82 9.0005
R5829 iovss.n107 iovss.n82 9.0005
R5830 iovss.n141 iovss.n82 9.0005
R5831 iovss.n106 iovss.n82 9.0005
R5832 iovss.n143 iovss.n82 9.0005
R5833 iovss.n105 iovss.n82 9.0005
R5834 iovss.n145 iovss.n82 9.0005
R5835 iovss.n104 iovss.n82 9.0005
R5836 iovss.n147 iovss.n82 9.0005
R5837 iovss.n82 iovss.n78 9.0005
R5838 iovss.n3436 iovss.n82 9.0005
R5839 iovss.n103 iovss.n82 9.0005
R5840 iovss.n3434 iovss.n82 9.0005
R5841 iovss.n82 iovss.n68 9.0005
R5842 iovss.n120 iovss.n91 9.0005
R5843 iovss.n118 iovss.n91 9.0005
R5844 iovss.n122 iovss.n91 9.0005
R5845 iovss.n117 iovss.n91 9.0005
R5846 iovss.n124 iovss.n91 9.0005
R5847 iovss.n116 iovss.n91 9.0005
R5848 iovss.n126 iovss.n91 9.0005
R5849 iovss.n115 iovss.n91 9.0005
R5850 iovss.n128 iovss.n91 9.0005
R5851 iovss.n114 iovss.n91 9.0005
R5852 iovss.n130 iovss.n91 9.0005
R5853 iovss.n113 iovss.n91 9.0005
R5854 iovss.n132 iovss.n91 9.0005
R5855 iovss.n112 iovss.n91 9.0005
R5856 iovss.n134 iovss.n91 9.0005
R5857 iovss.n111 iovss.n91 9.0005
R5858 iovss.n135 iovss.n91 9.0005
R5859 iovss.n110 iovss.n91 9.0005
R5860 iovss.n137 iovss.n91 9.0005
R5861 iovss.n109 iovss.n91 9.0005
R5862 iovss.n138 iovss.n91 9.0005
R5863 iovss.n108 iovss.n91 9.0005
R5864 iovss.n140 iovss.n91 9.0005
R5865 iovss.n107 iovss.n91 9.0005
R5866 iovss.n141 iovss.n91 9.0005
R5867 iovss.n106 iovss.n91 9.0005
R5868 iovss.n143 iovss.n91 9.0005
R5869 iovss.n105 iovss.n91 9.0005
R5870 iovss.n145 iovss.n91 9.0005
R5871 iovss.n104 iovss.n91 9.0005
R5872 iovss.n147 iovss.n91 9.0005
R5873 iovss.n91 iovss.n78 9.0005
R5874 iovss.n3436 iovss.n91 9.0005
R5875 iovss.n103 iovss.n91 9.0005
R5876 iovss.n3434 iovss.n91 9.0005
R5877 iovss.n91 iovss.n68 9.0005
R5878 iovss.n120 iovss.n81 9.0005
R5879 iovss.n118 iovss.n81 9.0005
R5880 iovss.n122 iovss.n81 9.0005
R5881 iovss.n117 iovss.n81 9.0005
R5882 iovss.n124 iovss.n81 9.0005
R5883 iovss.n116 iovss.n81 9.0005
R5884 iovss.n126 iovss.n81 9.0005
R5885 iovss.n115 iovss.n81 9.0005
R5886 iovss.n128 iovss.n81 9.0005
R5887 iovss.n114 iovss.n81 9.0005
R5888 iovss.n130 iovss.n81 9.0005
R5889 iovss.n113 iovss.n81 9.0005
R5890 iovss.n132 iovss.n81 9.0005
R5891 iovss.n112 iovss.n81 9.0005
R5892 iovss.n134 iovss.n81 9.0005
R5893 iovss.n111 iovss.n81 9.0005
R5894 iovss.n135 iovss.n81 9.0005
R5895 iovss.n110 iovss.n81 9.0005
R5896 iovss.n137 iovss.n81 9.0005
R5897 iovss.n109 iovss.n81 9.0005
R5898 iovss.n138 iovss.n81 9.0005
R5899 iovss.n108 iovss.n81 9.0005
R5900 iovss.n140 iovss.n81 9.0005
R5901 iovss.n107 iovss.n81 9.0005
R5902 iovss.n141 iovss.n81 9.0005
R5903 iovss.n106 iovss.n81 9.0005
R5904 iovss.n143 iovss.n81 9.0005
R5905 iovss.n105 iovss.n81 9.0005
R5906 iovss.n145 iovss.n81 9.0005
R5907 iovss.n104 iovss.n81 9.0005
R5908 iovss.n147 iovss.n81 9.0005
R5909 iovss.n81 iovss.n78 9.0005
R5910 iovss.n3436 iovss.n81 9.0005
R5911 iovss.n103 iovss.n81 9.0005
R5912 iovss.n3434 iovss.n81 9.0005
R5913 iovss.n81 iovss.n68 9.0005
R5914 iovss.n120 iovss.n92 9.0005
R5915 iovss.n118 iovss.n92 9.0005
R5916 iovss.n122 iovss.n92 9.0005
R5917 iovss.n117 iovss.n92 9.0005
R5918 iovss.n124 iovss.n92 9.0005
R5919 iovss.n116 iovss.n92 9.0005
R5920 iovss.n126 iovss.n92 9.0005
R5921 iovss.n115 iovss.n92 9.0005
R5922 iovss.n128 iovss.n92 9.0005
R5923 iovss.n114 iovss.n92 9.0005
R5924 iovss.n130 iovss.n92 9.0005
R5925 iovss.n113 iovss.n92 9.0005
R5926 iovss.n132 iovss.n92 9.0005
R5927 iovss.n112 iovss.n92 9.0005
R5928 iovss.n134 iovss.n92 9.0005
R5929 iovss.n111 iovss.n92 9.0005
R5930 iovss.n135 iovss.n92 9.0005
R5931 iovss.n110 iovss.n92 9.0005
R5932 iovss.n137 iovss.n92 9.0005
R5933 iovss.n109 iovss.n92 9.0005
R5934 iovss.n138 iovss.n92 9.0005
R5935 iovss.n108 iovss.n92 9.0005
R5936 iovss.n140 iovss.n92 9.0005
R5937 iovss.n107 iovss.n92 9.0005
R5938 iovss.n141 iovss.n92 9.0005
R5939 iovss.n106 iovss.n92 9.0005
R5940 iovss.n143 iovss.n92 9.0005
R5941 iovss.n105 iovss.n92 9.0005
R5942 iovss.n145 iovss.n92 9.0005
R5943 iovss.n104 iovss.n92 9.0005
R5944 iovss.n147 iovss.n92 9.0005
R5945 iovss.n92 iovss.n78 9.0005
R5946 iovss.n3436 iovss.n92 9.0005
R5947 iovss.n103 iovss.n92 9.0005
R5948 iovss.n3434 iovss.n92 9.0005
R5949 iovss.n92 iovss.n68 9.0005
R5950 iovss.n120 iovss.n80 9.0005
R5951 iovss.n118 iovss.n80 9.0005
R5952 iovss.n122 iovss.n80 9.0005
R5953 iovss.n117 iovss.n80 9.0005
R5954 iovss.n124 iovss.n80 9.0005
R5955 iovss.n116 iovss.n80 9.0005
R5956 iovss.n126 iovss.n80 9.0005
R5957 iovss.n115 iovss.n80 9.0005
R5958 iovss.n128 iovss.n80 9.0005
R5959 iovss.n114 iovss.n80 9.0005
R5960 iovss.n130 iovss.n80 9.0005
R5961 iovss.n113 iovss.n80 9.0005
R5962 iovss.n132 iovss.n80 9.0005
R5963 iovss.n112 iovss.n80 9.0005
R5964 iovss.n134 iovss.n80 9.0005
R5965 iovss.n111 iovss.n80 9.0005
R5966 iovss.n135 iovss.n80 9.0005
R5967 iovss.n110 iovss.n80 9.0005
R5968 iovss.n137 iovss.n80 9.0005
R5969 iovss.n109 iovss.n80 9.0005
R5970 iovss.n138 iovss.n80 9.0005
R5971 iovss.n108 iovss.n80 9.0005
R5972 iovss.n140 iovss.n80 9.0005
R5973 iovss.n107 iovss.n80 9.0005
R5974 iovss.n141 iovss.n80 9.0005
R5975 iovss.n106 iovss.n80 9.0005
R5976 iovss.n143 iovss.n80 9.0005
R5977 iovss.n105 iovss.n80 9.0005
R5978 iovss.n145 iovss.n80 9.0005
R5979 iovss.n104 iovss.n80 9.0005
R5980 iovss.n147 iovss.n80 9.0005
R5981 iovss.n80 iovss.n78 9.0005
R5982 iovss.n3436 iovss.n80 9.0005
R5983 iovss.n103 iovss.n80 9.0005
R5984 iovss.n3434 iovss.n80 9.0005
R5985 iovss.n80 iovss.n68 9.0005
R5986 iovss.n120 iovss.n93 9.0005
R5987 iovss.n118 iovss.n93 9.0005
R5988 iovss.n122 iovss.n93 9.0005
R5989 iovss.n117 iovss.n93 9.0005
R5990 iovss.n124 iovss.n93 9.0005
R5991 iovss.n116 iovss.n93 9.0005
R5992 iovss.n126 iovss.n93 9.0005
R5993 iovss.n115 iovss.n93 9.0005
R5994 iovss.n128 iovss.n93 9.0005
R5995 iovss.n114 iovss.n93 9.0005
R5996 iovss.n130 iovss.n93 9.0005
R5997 iovss.n113 iovss.n93 9.0005
R5998 iovss.n132 iovss.n93 9.0005
R5999 iovss.n112 iovss.n93 9.0005
R6000 iovss.n134 iovss.n93 9.0005
R6001 iovss.n111 iovss.n93 9.0005
R6002 iovss.n135 iovss.n93 9.0005
R6003 iovss.n110 iovss.n93 9.0005
R6004 iovss.n137 iovss.n93 9.0005
R6005 iovss.n109 iovss.n93 9.0005
R6006 iovss.n138 iovss.n93 9.0005
R6007 iovss.n108 iovss.n93 9.0005
R6008 iovss.n140 iovss.n93 9.0005
R6009 iovss.n107 iovss.n93 9.0005
R6010 iovss.n141 iovss.n93 9.0005
R6011 iovss.n106 iovss.n93 9.0005
R6012 iovss.n143 iovss.n93 9.0005
R6013 iovss.n105 iovss.n93 9.0005
R6014 iovss.n145 iovss.n93 9.0005
R6015 iovss.n104 iovss.n93 9.0005
R6016 iovss.n147 iovss.n93 9.0005
R6017 iovss.n93 iovss.n78 9.0005
R6018 iovss.n3436 iovss.n93 9.0005
R6019 iovss.n103 iovss.n93 9.0005
R6020 iovss.n3434 iovss.n93 9.0005
R6021 iovss.n93 iovss.n68 9.0005
R6022 iovss.n120 iovss.n79 9.0005
R6023 iovss.n118 iovss.n79 9.0005
R6024 iovss.n122 iovss.n79 9.0005
R6025 iovss.n117 iovss.n79 9.0005
R6026 iovss.n124 iovss.n79 9.0005
R6027 iovss.n116 iovss.n79 9.0005
R6028 iovss.n126 iovss.n79 9.0005
R6029 iovss.n115 iovss.n79 9.0005
R6030 iovss.n128 iovss.n79 9.0005
R6031 iovss.n114 iovss.n79 9.0005
R6032 iovss.n130 iovss.n79 9.0005
R6033 iovss.n113 iovss.n79 9.0005
R6034 iovss.n132 iovss.n79 9.0005
R6035 iovss.n112 iovss.n79 9.0005
R6036 iovss.n134 iovss.n79 9.0005
R6037 iovss.n111 iovss.n79 9.0005
R6038 iovss.n135 iovss.n79 9.0005
R6039 iovss.n110 iovss.n79 9.0005
R6040 iovss.n137 iovss.n79 9.0005
R6041 iovss.n109 iovss.n79 9.0005
R6042 iovss.n138 iovss.n79 9.0005
R6043 iovss.n108 iovss.n79 9.0005
R6044 iovss.n140 iovss.n79 9.0005
R6045 iovss.n107 iovss.n79 9.0005
R6046 iovss.n141 iovss.n79 9.0005
R6047 iovss.n106 iovss.n79 9.0005
R6048 iovss.n143 iovss.n79 9.0005
R6049 iovss.n105 iovss.n79 9.0005
R6050 iovss.n145 iovss.n79 9.0005
R6051 iovss.n104 iovss.n79 9.0005
R6052 iovss.n147 iovss.n79 9.0005
R6053 iovss.n79 iovss.n78 9.0005
R6054 iovss.n3436 iovss.n79 9.0005
R6055 iovss.n103 iovss.n79 9.0005
R6056 iovss.n3434 iovss.n79 9.0005
R6057 iovss.n79 iovss.n68 9.0005
R6058 iovss.n3435 iovss.n120 9.0005
R6059 iovss.n3435 iovss.n118 9.0005
R6060 iovss.n3435 iovss.n122 9.0005
R6061 iovss.n3435 iovss.n117 9.0005
R6062 iovss.n3435 iovss.n124 9.0005
R6063 iovss.n3435 iovss.n116 9.0005
R6064 iovss.n3435 iovss.n126 9.0005
R6065 iovss.n3435 iovss.n115 9.0005
R6066 iovss.n3435 iovss.n128 9.0005
R6067 iovss.n3435 iovss.n114 9.0005
R6068 iovss.n3435 iovss.n130 9.0005
R6069 iovss.n3435 iovss.n113 9.0005
R6070 iovss.n3435 iovss.n132 9.0005
R6071 iovss.n3435 iovss.n112 9.0005
R6072 iovss.n3435 iovss.n134 9.0005
R6073 iovss.n3435 iovss.n111 9.0005
R6074 iovss.n3435 iovss.n135 9.0005
R6075 iovss.n3435 iovss.n110 9.0005
R6076 iovss.n3435 iovss.n137 9.0005
R6077 iovss.n3435 iovss.n109 9.0005
R6078 iovss.n3435 iovss.n138 9.0005
R6079 iovss.n3435 iovss.n108 9.0005
R6080 iovss.n3435 iovss.n140 9.0005
R6081 iovss.n3435 iovss.n107 9.0005
R6082 iovss.n3435 iovss.n141 9.0005
R6083 iovss.n3435 iovss.n106 9.0005
R6084 iovss.n3435 iovss.n143 9.0005
R6085 iovss.n3435 iovss.n105 9.0005
R6086 iovss.n3435 iovss.n145 9.0005
R6087 iovss.n3435 iovss.n104 9.0005
R6088 iovss.n3435 iovss.n147 9.0005
R6089 iovss.n3435 iovss.n78 9.0005
R6090 iovss.n3436 iovss.n3435 9.0005
R6091 iovss.n3435 iovss.n103 9.0005
R6092 iovss.n3435 iovss.n3434 9.0005
R6093 iovss.n3435 iovss.n101 9.0005
R6094 iovss.n3435 iovss.n68 9.0005
R6095 iovss.n1596 iovss.n220 9.0005
R6096 iovss.n1553 iovss.n220 9.0005
R6097 iovss.n1599 iovss.n220 9.0005
R6098 iovss.n1551 iovss.n220 9.0005
R6099 iovss.n2394 iovss.n220 9.0005
R6100 iovss.n2393 iovss.n1569 9.0005
R6101 iovss.n2393 iovss.n1566 9.0005
R6102 iovss.n2393 iovss.n1573 9.0005
R6103 iovss.n2393 iovss.n1564 9.0005
R6104 iovss.n2393 iovss.n1577 9.0005
R6105 iovss.n2393 iovss.n1562 9.0005
R6106 iovss.n2393 iovss.n1581 9.0005
R6107 iovss.n2393 iovss.n1560 9.0005
R6108 iovss.n2393 iovss.n1585 9.0005
R6109 iovss.n2393 iovss.n1558 9.0005
R6110 iovss.n2393 iovss.n1589 9.0005
R6111 iovss.n2394 iovss.n2393 9.0005
R6112 iovss.n1624 iovss.n1569 9.0005
R6113 iovss.n1624 iovss.n1567 9.0005
R6114 iovss.n1624 iovss.n1571 9.0005
R6115 iovss.n1624 iovss.n1566 9.0005
R6116 iovss.n1624 iovss.n1573 9.0005
R6117 iovss.n1624 iovss.n1565 9.0005
R6118 iovss.n1624 iovss.n1575 9.0005
R6119 iovss.n1624 iovss.n1564 9.0005
R6120 iovss.n1624 iovss.n1577 9.0005
R6121 iovss.n1624 iovss.n1563 9.0005
R6122 iovss.n1624 iovss.n1579 9.0005
R6123 iovss.n1624 iovss.n1562 9.0005
R6124 iovss.n1624 iovss.n1581 9.0005
R6125 iovss.n1624 iovss.n1561 9.0005
R6126 iovss.n1624 iovss.n1583 9.0005
R6127 iovss.n1624 iovss.n1560 9.0005
R6128 iovss.n1624 iovss.n1585 9.0005
R6129 iovss.n1624 iovss.n1559 9.0005
R6130 iovss.n1624 iovss.n1587 9.0005
R6131 iovss.n1624 iovss.n1558 9.0005
R6132 iovss.n1624 iovss.n1589 9.0005
R6133 iovss.n1624 iovss.n1557 9.0005
R6134 iovss.n1624 iovss.n1591 9.0005
R6135 iovss.n1624 iovss.n1556 9.0005
R6136 iovss.n1624 iovss.n1593 9.0005
R6137 iovss.n1624 iovss.n1555 9.0005
R6138 iovss.n1624 iovss.n1595 9.0005
R6139 iovss.n1624 iovss.n1554 9.0005
R6140 iovss.n1624 iovss.n1596 9.0005
R6141 iovss.n1624 iovss.n1553 9.0005
R6142 iovss.n1624 iovss.n1598 9.0005
R6143 iovss.n1624 iovss.n1552 9.0005
R6144 iovss.n1624 iovss.n1599 9.0005
R6145 iovss.n1624 iovss.n1551 9.0005
R6146 iovss.n2396 iovss.n1624 9.0005
R6147 iovss.n2394 iovss.n1624 9.0005
R6148 iovss.n1627 iovss.n1569 9.0005
R6149 iovss.n1627 iovss.n1567 9.0005
R6150 iovss.n1627 iovss.n1571 9.0005
R6151 iovss.n1627 iovss.n1566 9.0005
R6152 iovss.n1627 iovss.n1573 9.0005
R6153 iovss.n1627 iovss.n1565 9.0005
R6154 iovss.n1627 iovss.n1575 9.0005
R6155 iovss.n1627 iovss.n1564 9.0005
R6156 iovss.n1627 iovss.n1577 9.0005
R6157 iovss.n1627 iovss.n1563 9.0005
R6158 iovss.n1627 iovss.n1579 9.0005
R6159 iovss.n1627 iovss.n1562 9.0005
R6160 iovss.n1627 iovss.n1581 9.0005
R6161 iovss.n1627 iovss.n1561 9.0005
R6162 iovss.n1627 iovss.n1583 9.0005
R6163 iovss.n1627 iovss.n1560 9.0005
R6164 iovss.n1627 iovss.n1585 9.0005
R6165 iovss.n1627 iovss.n1559 9.0005
R6166 iovss.n1627 iovss.n1587 9.0005
R6167 iovss.n1627 iovss.n1558 9.0005
R6168 iovss.n1627 iovss.n1589 9.0005
R6169 iovss.n1627 iovss.n1557 9.0005
R6170 iovss.n1627 iovss.n1591 9.0005
R6171 iovss.n1627 iovss.n1556 9.0005
R6172 iovss.n1627 iovss.n1593 9.0005
R6173 iovss.n1627 iovss.n1555 9.0005
R6174 iovss.n1627 iovss.n1595 9.0005
R6175 iovss.n1627 iovss.n1554 9.0005
R6176 iovss.n1627 iovss.n1596 9.0005
R6177 iovss.n1627 iovss.n1553 9.0005
R6178 iovss.n1627 iovss.n1598 9.0005
R6179 iovss.n1627 iovss.n1552 9.0005
R6180 iovss.n1627 iovss.n1599 9.0005
R6181 iovss.n1627 iovss.n1551 9.0005
R6182 iovss.n2396 iovss.n1627 9.0005
R6183 iovss.n2394 iovss.n1627 9.0005
R6184 iovss.n1623 iovss.n1569 9.0005
R6185 iovss.n1623 iovss.n1567 9.0005
R6186 iovss.n1623 iovss.n1571 9.0005
R6187 iovss.n1623 iovss.n1566 9.0005
R6188 iovss.n1623 iovss.n1573 9.0005
R6189 iovss.n1623 iovss.n1565 9.0005
R6190 iovss.n1623 iovss.n1575 9.0005
R6191 iovss.n1623 iovss.n1564 9.0005
R6192 iovss.n1623 iovss.n1577 9.0005
R6193 iovss.n1623 iovss.n1563 9.0005
R6194 iovss.n1623 iovss.n1579 9.0005
R6195 iovss.n1623 iovss.n1562 9.0005
R6196 iovss.n1623 iovss.n1581 9.0005
R6197 iovss.n1623 iovss.n1561 9.0005
R6198 iovss.n1623 iovss.n1583 9.0005
R6199 iovss.n1623 iovss.n1560 9.0005
R6200 iovss.n1623 iovss.n1585 9.0005
R6201 iovss.n1623 iovss.n1559 9.0005
R6202 iovss.n1623 iovss.n1587 9.0005
R6203 iovss.n1623 iovss.n1558 9.0005
R6204 iovss.n1623 iovss.n1589 9.0005
R6205 iovss.n1623 iovss.n1557 9.0005
R6206 iovss.n1623 iovss.n1591 9.0005
R6207 iovss.n1623 iovss.n1556 9.0005
R6208 iovss.n1623 iovss.n1593 9.0005
R6209 iovss.n1623 iovss.n1555 9.0005
R6210 iovss.n1623 iovss.n1595 9.0005
R6211 iovss.n1623 iovss.n1554 9.0005
R6212 iovss.n1623 iovss.n1596 9.0005
R6213 iovss.n1623 iovss.n1553 9.0005
R6214 iovss.n1623 iovss.n1598 9.0005
R6215 iovss.n1623 iovss.n1552 9.0005
R6216 iovss.n1623 iovss.n1599 9.0005
R6217 iovss.n1623 iovss.n1551 9.0005
R6218 iovss.n2396 iovss.n1623 9.0005
R6219 iovss.n2394 iovss.n1623 9.0005
R6220 iovss.n1628 iovss.n1569 9.0005
R6221 iovss.n1628 iovss.n1567 9.0005
R6222 iovss.n1628 iovss.n1571 9.0005
R6223 iovss.n1628 iovss.n1566 9.0005
R6224 iovss.n1628 iovss.n1573 9.0005
R6225 iovss.n1628 iovss.n1565 9.0005
R6226 iovss.n1628 iovss.n1575 9.0005
R6227 iovss.n1628 iovss.n1564 9.0005
R6228 iovss.n1628 iovss.n1577 9.0005
R6229 iovss.n1628 iovss.n1563 9.0005
R6230 iovss.n1628 iovss.n1579 9.0005
R6231 iovss.n1628 iovss.n1562 9.0005
R6232 iovss.n1628 iovss.n1581 9.0005
R6233 iovss.n1628 iovss.n1561 9.0005
R6234 iovss.n1628 iovss.n1583 9.0005
R6235 iovss.n1628 iovss.n1560 9.0005
R6236 iovss.n1628 iovss.n1585 9.0005
R6237 iovss.n1628 iovss.n1559 9.0005
R6238 iovss.n1628 iovss.n1587 9.0005
R6239 iovss.n1628 iovss.n1558 9.0005
R6240 iovss.n1628 iovss.n1589 9.0005
R6241 iovss.n1628 iovss.n1557 9.0005
R6242 iovss.n1628 iovss.n1591 9.0005
R6243 iovss.n1628 iovss.n1556 9.0005
R6244 iovss.n1628 iovss.n1593 9.0005
R6245 iovss.n1628 iovss.n1555 9.0005
R6246 iovss.n1628 iovss.n1595 9.0005
R6247 iovss.n1628 iovss.n1554 9.0005
R6248 iovss.n1628 iovss.n1596 9.0005
R6249 iovss.n1628 iovss.n1553 9.0005
R6250 iovss.n1628 iovss.n1598 9.0005
R6251 iovss.n1628 iovss.n1552 9.0005
R6252 iovss.n1628 iovss.n1599 9.0005
R6253 iovss.n1628 iovss.n1551 9.0005
R6254 iovss.n2396 iovss.n1628 9.0005
R6255 iovss.n2394 iovss.n1628 9.0005
R6256 iovss.n1622 iovss.n1569 9.0005
R6257 iovss.n1622 iovss.n1567 9.0005
R6258 iovss.n1622 iovss.n1571 9.0005
R6259 iovss.n1622 iovss.n1566 9.0005
R6260 iovss.n1622 iovss.n1573 9.0005
R6261 iovss.n1622 iovss.n1565 9.0005
R6262 iovss.n1622 iovss.n1575 9.0005
R6263 iovss.n1622 iovss.n1564 9.0005
R6264 iovss.n1622 iovss.n1577 9.0005
R6265 iovss.n1622 iovss.n1563 9.0005
R6266 iovss.n1622 iovss.n1579 9.0005
R6267 iovss.n1622 iovss.n1562 9.0005
R6268 iovss.n1622 iovss.n1581 9.0005
R6269 iovss.n1622 iovss.n1561 9.0005
R6270 iovss.n1622 iovss.n1583 9.0005
R6271 iovss.n1622 iovss.n1560 9.0005
R6272 iovss.n1622 iovss.n1585 9.0005
R6273 iovss.n1622 iovss.n1559 9.0005
R6274 iovss.n1622 iovss.n1587 9.0005
R6275 iovss.n1622 iovss.n1558 9.0005
R6276 iovss.n1622 iovss.n1589 9.0005
R6277 iovss.n1622 iovss.n1557 9.0005
R6278 iovss.n1622 iovss.n1591 9.0005
R6279 iovss.n1622 iovss.n1556 9.0005
R6280 iovss.n1622 iovss.n1593 9.0005
R6281 iovss.n1622 iovss.n1555 9.0005
R6282 iovss.n1622 iovss.n1595 9.0005
R6283 iovss.n1622 iovss.n1554 9.0005
R6284 iovss.n1622 iovss.n1596 9.0005
R6285 iovss.n1622 iovss.n1553 9.0005
R6286 iovss.n1622 iovss.n1598 9.0005
R6287 iovss.n1622 iovss.n1552 9.0005
R6288 iovss.n1622 iovss.n1599 9.0005
R6289 iovss.n1622 iovss.n1551 9.0005
R6290 iovss.n2396 iovss.n1622 9.0005
R6291 iovss.n2394 iovss.n1622 9.0005
R6292 iovss.n1629 iovss.n1569 9.0005
R6293 iovss.n1629 iovss.n1567 9.0005
R6294 iovss.n1629 iovss.n1571 9.0005
R6295 iovss.n1629 iovss.n1566 9.0005
R6296 iovss.n1629 iovss.n1573 9.0005
R6297 iovss.n1629 iovss.n1565 9.0005
R6298 iovss.n1629 iovss.n1575 9.0005
R6299 iovss.n1629 iovss.n1564 9.0005
R6300 iovss.n1629 iovss.n1577 9.0005
R6301 iovss.n1629 iovss.n1563 9.0005
R6302 iovss.n1629 iovss.n1579 9.0005
R6303 iovss.n1629 iovss.n1562 9.0005
R6304 iovss.n1629 iovss.n1581 9.0005
R6305 iovss.n1629 iovss.n1561 9.0005
R6306 iovss.n1629 iovss.n1583 9.0005
R6307 iovss.n1629 iovss.n1560 9.0005
R6308 iovss.n1629 iovss.n1585 9.0005
R6309 iovss.n1629 iovss.n1559 9.0005
R6310 iovss.n1629 iovss.n1587 9.0005
R6311 iovss.n1629 iovss.n1558 9.0005
R6312 iovss.n1629 iovss.n1589 9.0005
R6313 iovss.n1629 iovss.n1557 9.0005
R6314 iovss.n1629 iovss.n1591 9.0005
R6315 iovss.n1629 iovss.n1556 9.0005
R6316 iovss.n1629 iovss.n1593 9.0005
R6317 iovss.n1629 iovss.n1555 9.0005
R6318 iovss.n1629 iovss.n1595 9.0005
R6319 iovss.n1629 iovss.n1554 9.0005
R6320 iovss.n1629 iovss.n1596 9.0005
R6321 iovss.n1629 iovss.n1553 9.0005
R6322 iovss.n1629 iovss.n1598 9.0005
R6323 iovss.n1629 iovss.n1552 9.0005
R6324 iovss.n1629 iovss.n1599 9.0005
R6325 iovss.n1629 iovss.n1551 9.0005
R6326 iovss.n2396 iovss.n1629 9.0005
R6327 iovss.n2394 iovss.n1629 9.0005
R6328 iovss.n1621 iovss.n1569 9.0005
R6329 iovss.n1621 iovss.n1567 9.0005
R6330 iovss.n1621 iovss.n1571 9.0005
R6331 iovss.n1621 iovss.n1566 9.0005
R6332 iovss.n1621 iovss.n1573 9.0005
R6333 iovss.n1621 iovss.n1565 9.0005
R6334 iovss.n1621 iovss.n1575 9.0005
R6335 iovss.n1621 iovss.n1564 9.0005
R6336 iovss.n1621 iovss.n1577 9.0005
R6337 iovss.n1621 iovss.n1563 9.0005
R6338 iovss.n1621 iovss.n1579 9.0005
R6339 iovss.n1621 iovss.n1562 9.0005
R6340 iovss.n1621 iovss.n1581 9.0005
R6341 iovss.n1621 iovss.n1561 9.0005
R6342 iovss.n1621 iovss.n1583 9.0005
R6343 iovss.n1621 iovss.n1560 9.0005
R6344 iovss.n1621 iovss.n1585 9.0005
R6345 iovss.n1621 iovss.n1559 9.0005
R6346 iovss.n1621 iovss.n1587 9.0005
R6347 iovss.n1621 iovss.n1558 9.0005
R6348 iovss.n1621 iovss.n1589 9.0005
R6349 iovss.n1621 iovss.n1557 9.0005
R6350 iovss.n1621 iovss.n1591 9.0005
R6351 iovss.n1621 iovss.n1556 9.0005
R6352 iovss.n1621 iovss.n1593 9.0005
R6353 iovss.n1621 iovss.n1555 9.0005
R6354 iovss.n1621 iovss.n1595 9.0005
R6355 iovss.n1621 iovss.n1554 9.0005
R6356 iovss.n1621 iovss.n1596 9.0005
R6357 iovss.n1621 iovss.n1553 9.0005
R6358 iovss.n1621 iovss.n1598 9.0005
R6359 iovss.n1621 iovss.n1552 9.0005
R6360 iovss.n1621 iovss.n1599 9.0005
R6361 iovss.n1621 iovss.n1551 9.0005
R6362 iovss.n2396 iovss.n1621 9.0005
R6363 iovss.n2394 iovss.n1621 9.0005
R6364 iovss.n1630 iovss.n1569 9.0005
R6365 iovss.n1630 iovss.n1567 9.0005
R6366 iovss.n1630 iovss.n1571 9.0005
R6367 iovss.n1630 iovss.n1566 9.0005
R6368 iovss.n1630 iovss.n1573 9.0005
R6369 iovss.n1630 iovss.n1565 9.0005
R6370 iovss.n1630 iovss.n1575 9.0005
R6371 iovss.n1630 iovss.n1564 9.0005
R6372 iovss.n1630 iovss.n1577 9.0005
R6373 iovss.n1630 iovss.n1563 9.0005
R6374 iovss.n1630 iovss.n1579 9.0005
R6375 iovss.n1630 iovss.n1562 9.0005
R6376 iovss.n1630 iovss.n1581 9.0005
R6377 iovss.n1630 iovss.n1561 9.0005
R6378 iovss.n1630 iovss.n1583 9.0005
R6379 iovss.n1630 iovss.n1560 9.0005
R6380 iovss.n1630 iovss.n1585 9.0005
R6381 iovss.n1630 iovss.n1559 9.0005
R6382 iovss.n1630 iovss.n1587 9.0005
R6383 iovss.n1630 iovss.n1558 9.0005
R6384 iovss.n1630 iovss.n1589 9.0005
R6385 iovss.n1630 iovss.n1557 9.0005
R6386 iovss.n1630 iovss.n1591 9.0005
R6387 iovss.n1630 iovss.n1556 9.0005
R6388 iovss.n1630 iovss.n1593 9.0005
R6389 iovss.n1630 iovss.n1555 9.0005
R6390 iovss.n1630 iovss.n1595 9.0005
R6391 iovss.n1630 iovss.n1554 9.0005
R6392 iovss.n1630 iovss.n1596 9.0005
R6393 iovss.n1630 iovss.n1553 9.0005
R6394 iovss.n1630 iovss.n1598 9.0005
R6395 iovss.n1630 iovss.n1552 9.0005
R6396 iovss.n1630 iovss.n1599 9.0005
R6397 iovss.n1630 iovss.n1551 9.0005
R6398 iovss.n2396 iovss.n1630 9.0005
R6399 iovss.n2394 iovss.n1630 9.0005
R6400 iovss.n1620 iovss.n1569 9.0005
R6401 iovss.n1620 iovss.n1567 9.0005
R6402 iovss.n1620 iovss.n1571 9.0005
R6403 iovss.n1620 iovss.n1566 9.0005
R6404 iovss.n1620 iovss.n1573 9.0005
R6405 iovss.n1620 iovss.n1565 9.0005
R6406 iovss.n1620 iovss.n1575 9.0005
R6407 iovss.n1620 iovss.n1564 9.0005
R6408 iovss.n1620 iovss.n1577 9.0005
R6409 iovss.n1620 iovss.n1563 9.0005
R6410 iovss.n1620 iovss.n1579 9.0005
R6411 iovss.n1620 iovss.n1562 9.0005
R6412 iovss.n1620 iovss.n1581 9.0005
R6413 iovss.n1620 iovss.n1561 9.0005
R6414 iovss.n1620 iovss.n1583 9.0005
R6415 iovss.n1620 iovss.n1560 9.0005
R6416 iovss.n1620 iovss.n1585 9.0005
R6417 iovss.n1620 iovss.n1559 9.0005
R6418 iovss.n1620 iovss.n1587 9.0005
R6419 iovss.n1620 iovss.n1558 9.0005
R6420 iovss.n1620 iovss.n1589 9.0005
R6421 iovss.n1620 iovss.n1557 9.0005
R6422 iovss.n1620 iovss.n1591 9.0005
R6423 iovss.n1620 iovss.n1556 9.0005
R6424 iovss.n1620 iovss.n1593 9.0005
R6425 iovss.n1620 iovss.n1555 9.0005
R6426 iovss.n1620 iovss.n1595 9.0005
R6427 iovss.n1620 iovss.n1554 9.0005
R6428 iovss.n1620 iovss.n1596 9.0005
R6429 iovss.n1620 iovss.n1553 9.0005
R6430 iovss.n1620 iovss.n1598 9.0005
R6431 iovss.n1620 iovss.n1552 9.0005
R6432 iovss.n1620 iovss.n1599 9.0005
R6433 iovss.n1620 iovss.n1551 9.0005
R6434 iovss.n2396 iovss.n1620 9.0005
R6435 iovss.n2394 iovss.n1620 9.0005
R6436 iovss.n1631 iovss.n1569 9.0005
R6437 iovss.n1631 iovss.n1567 9.0005
R6438 iovss.n1631 iovss.n1571 9.0005
R6439 iovss.n1631 iovss.n1566 9.0005
R6440 iovss.n1631 iovss.n1573 9.0005
R6441 iovss.n1631 iovss.n1565 9.0005
R6442 iovss.n1631 iovss.n1575 9.0005
R6443 iovss.n1631 iovss.n1564 9.0005
R6444 iovss.n1631 iovss.n1577 9.0005
R6445 iovss.n1631 iovss.n1563 9.0005
R6446 iovss.n1631 iovss.n1579 9.0005
R6447 iovss.n1631 iovss.n1562 9.0005
R6448 iovss.n1631 iovss.n1581 9.0005
R6449 iovss.n1631 iovss.n1561 9.0005
R6450 iovss.n1631 iovss.n1583 9.0005
R6451 iovss.n1631 iovss.n1560 9.0005
R6452 iovss.n1631 iovss.n1585 9.0005
R6453 iovss.n1631 iovss.n1559 9.0005
R6454 iovss.n1631 iovss.n1587 9.0005
R6455 iovss.n1631 iovss.n1558 9.0005
R6456 iovss.n1631 iovss.n1589 9.0005
R6457 iovss.n1631 iovss.n1557 9.0005
R6458 iovss.n1631 iovss.n1591 9.0005
R6459 iovss.n1631 iovss.n1556 9.0005
R6460 iovss.n1631 iovss.n1593 9.0005
R6461 iovss.n1631 iovss.n1555 9.0005
R6462 iovss.n1631 iovss.n1595 9.0005
R6463 iovss.n1631 iovss.n1554 9.0005
R6464 iovss.n1631 iovss.n1596 9.0005
R6465 iovss.n1631 iovss.n1553 9.0005
R6466 iovss.n1631 iovss.n1598 9.0005
R6467 iovss.n1631 iovss.n1552 9.0005
R6468 iovss.n1631 iovss.n1599 9.0005
R6469 iovss.n1631 iovss.n1551 9.0005
R6470 iovss.n2396 iovss.n1631 9.0005
R6471 iovss.n2394 iovss.n1631 9.0005
R6472 iovss.n1619 iovss.n1569 9.0005
R6473 iovss.n1619 iovss.n1567 9.0005
R6474 iovss.n1619 iovss.n1571 9.0005
R6475 iovss.n1619 iovss.n1566 9.0005
R6476 iovss.n1619 iovss.n1573 9.0005
R6477 iovss.n1619 iovss.n1565 9.0005
R6478 iovss.n1619 iovss.n1575 9.0005
R6479 iovss.n1619 iovss.n1564 9.0005
R6480 iovss.n1619 iovss.n1577 9.0005
R6481 iovss.n1619 iovss.n1563 9.0005
R6482 iovss.n1619 iovss.n1579 9.0005
R6483 iovss.n1619 iovss.n1562 9.0005
R6484 iovss.n1619 iovss.n1581 9.0005
R6485 iovss.n1619 iovss.n1561 9.0005
R6486 iovss.n1619 iovss.n1583 9.0005
R6487 iovss.n1619 iovss.n1560 9.0005
R6488 iovss.n1619 iovss.n1585 9.0005
R6489 iovss.n1619 iovss.n1559 9.0005
R6490 iovss.n1619 iovss.n1587 9.0005
R6491 iovss.n1619 iovss.n1558 9.0005
R6492 iovss.n1619 iovss.n1589 9.0005
R6493 iovss.n1619 iovss.n1557 9.0005
R6494 iovss.n1619 iovss.n1591 9.0005
R6495 iovss.n1619 iovss.n1556 9.0005
R6496 iovss.n1619 iovss.n1593 9.0005
R6497 iovss.n1619 iovss.n1555 9.0005
R6498 iovss.n1619 iovss.n1595 9.0005
R6499 iovss.n1619 iovss.n1554 9.0005
R6500 iovss.n1619 iovss.n1596 9.0005
R6501 iovss.n1619 iovss.n1553 9.0005
R6502 iovss.n1619 iovss.n1598 9.0005
R6503 iovss.n1619 iovss.n1552 9.0005
R6504 iovss.n1619 iovss.n1599 9.0005
R6505 iovss.n1619 iovss.n1551 9.0005
R6506 iovss.n2396 iovss.n1619 9.0005
R6507 iovss.n2394 iovss.n1619 9.0005
R6508 iovss.n1632 iovss.n1569 9.0005
R6509 iovss.n1632 iovss.n1567 9.0005
R6510 iovss.n1632 iovss.n1571 9.0005
R6511 iovss.n1632 iovss.n1566 9.0005
R6512 iovss.n1632 iovss.n1573 9.0005
R6513 iovss.n1632 iovss.n1565 9.0005
R6514 iovss.n1632 iovss.n1575 9.0005
R6515 iovss.n1632 iovss.n1564 9.0005
R6516 iovss.n1632 iovss.n1577 9.0005
R6517 iovss.n1632 iovss.n1563 9.0005
R6518 iovss.n1632 iovss.n1579 9.0005
R6519 iovss.n1632 iovss.n1562 9.0005
R6520 iovss.n1632 iovss.n1581 9.0005
R6521 iovss.n1632 iovss.n1561 9.0005
R6522 iovss.n1632 iovss.n1583 9.0005
R6523 iovss.n1632 iovss.n1560 9.0005
R6524 iovss.n1632 iovss.n1585 9.0005
R6525 iovss.n1632 iovss.n1559 9.0005
R6526 iovss.n1632 iovss.n1587 9.0005
R6527 iovss.n1632 iovss.n1558 9.0005
R6528 iovss.n1632 iovss.n1589 9.0005
R6529 iovss.n1632 iovss.n1557 9.0005
R6530 iovss.n1632 iovss.n1591 9.0005
R6531 iovss.n1632 iovss.n1556 9.0005
R6532 iovss.n1632 iovss.n1593 9.0005
R6533 iovss.n1632 iovss.n1555 9.0005
R6534 iovss.n1632 iovss.n1595 9.0005
R6535 iovss.n1632 iovss.n1554 9.0005
R6536 iovss.n1632 iovss.n1596 9.0005
R6537 iovss.n1632 iovss.n1553 9.0005
R6538 iovss.n1632 iovss.n1598 9.0005
R6539 iovss.n1632 iovss.n1552 9.0005
R6540 iovss.n1632 iovss.n1599 9.0005
R6541 iovss.n1632 iovss.n1551 9.0005
R6542 iovss.n2396 iovss.n1632 9.0005
R6543 iovss.n2394 iovss.n1632 9.0005
R6544 iovss.n1618 iovss.n1569 9.0005
R6545 iovss.n1618 iovss.n1567 9.0005
R6546 iovss.n1618 iovss.n1571 9.0005
R6547 iovss.n1618 iovss.n1566 9.0005
R6548 iovss.n1618 iovss.n1573 9.0005
R6549 iovss.n1618 iovss.n1565 9.0005
R6550 iovss.n1618 iovss.n1575 9.0005
R6551 iovss.n1618 iovss.n1564 9.0005
R6552 iovss.n1618 iovss.n1577 9.0005
R6553 iovss.n1618 iovss.n1563 9.0005
R6554 iovss.n1618 iovss.n1579 9.0005
R6555 iovss.n1618 iovss.n1562 9.0005
R6556 iovss.n1618 iovss.n1581 9.0005
R6557 iovss.n1618 iovss.n1561 9.0005
R6558 iovss.n1618 iovss.n1583 9.0005
R6559 iovss.n1618 iovss.n1560 9.0005
R6560 iovss.n1618 iovss.n1585 9.0005
R6561 iovss.n1618 iovss.n1559 9.0005
R6562 iovss.n1618 iovss.n1587 9.0005
R6563 iovss.n1618 iovss.n1558 9.0005
R6564 iovss.n1618 iovss.n1589 9.0005
R6565 iovss.n1618 iovss.n1557 9.0005
R6566 iovss.n1618 iovss.n1591 9.0005
R6567 iovss.n1618 iovss.n1556 9.0005
R6568 iovss.n1618 iovss.n1593 9.0005
R6569 iovss.n1618 iovss.n1555 9.0005
R6570 iovss.n1618 iovss.n1595 9.0005
R6571 iovss.n1618 iovss.n1554 9.0005
R6572 iovss.n1618 iovss.n1596 9.0005
R6573 iovss.n1618 iovss.n1553 9.0005
R6574 iovss.n1618 iovss.n1598 9.0005
R6575 iovss.n1618 iovss.n1552 9.0005
R6576 iovss.n1618 iovss.n1599 9.0005
R6577 iovss.n1618 iovss.n1551 9.0005
R6578 iovss.n2396 iovss.n1618 9.0005
R6579 iovss.n2394 iovss.n1618 9.0005
R6580 iovss.n1633 iovss.n1569 9.0005
R6581 iovss.n1633 iovss.n1567 9.0005
R6582 iovss.n1633 iovss.n1571 9.0005
R6583 iovss.n1633 iovss.n1566 9.0005
R6584 iovss.n1633 iovss.n1573 9.0005
R6585 iovss.n1633 iovss.n1565 9.0005
R6586 iovss.n1633 iovss.n1575 9.0005
R6587 iovss.n1633 iovss.n1564 9.0005
R6588 iovss.n1633 iovss.n1577 9.0005
R6589 iovss.n1633 iovss.n1563 9.0005
R6590 iovss.n1633 iovss.n1579 9.0005
R6591 iovss.n1633 iovss.n1562 9.0005
R6592 iovss.n1633 iovss.n1581 9.0005
R6593 iovss.n1633 iovss.n1561 9.0005
R6594 iovss.n1633 iovss.n1583 9.0005
R6595 iovss.n1633 iovss.n1560 9.0005
R6596 iovss.n1633 iovss.n1585 9.0005
R6597 iovss.n1633 iovss.n1559 9.0005
R6598 iovss.n1633 iovss.n1587 9.0005
R6599 iovss.n1633 iovss.n1558 9.0005
R6600 iovss.n1633 iovss.n1589 9.0005
R6601 iovss.n1633 iovss.n1557 9.0005
R6602 iovss.n1633 iovss.n1591 9.0005
R6603 iovss.n1633 iovss.n1556 9.0005
R6604 iovss.n1633 iovss.n1593 9.0005
R6605 iovss.n1633 iovss.n1555 9.0005
R6606 iovss.n1633 iovss.n1595 9.0005
R6607 iovss.n1633 iovss.n1554 9.0005
R6608 iovss.n1633 iovss.n1596 9.0005
R6609 iovss.n1633 iovss.n1553 9.0005
R6610 iovss.n1633 iovss.n1598 9.0005
R6611 iovss.n1633 iovss.n1552 9.0005
R6612 iovss.n1633 iovss.n1599 9.0005
R6613 iovss.n1633 iovss.n1551 9.0005
R6614 iovss.n2396 iovss.n1633 9.0005
R6615 iovss.n2394 iovss.n1633 9.0005
R6616 iovss.n1617 iovss.n1569 9.0005
R6617 iovss.n1617 iovss.n1567 9.0005
R6618 iovss.n1617 iovss.n1571 9.0005
R6619 iovss.n1617 iovss.n1566 9.0005
R6620 iovss.n1617 iovss.n1573 9.0005
R6621 iovss.n1617 iovss.n1565 9.0005
R6622 iovss.n1617 iovss.n1575 9.0005
R6623 iovss.n1617 iovss.n1564 9.0005
R6624 iovss.n1617 iovss.n1577 9.0005
R6625 iovss.n1617 iovss.n1563 9.0005
R6626 iovss.n1617 iovss.n1579 9.0005
R6627 iovss.n1617 iovss.n1562 9.0005
R6628 iovss.n1617 iovss.n1581 9.0005
R6629 iovss.n1617 iovss.n1561 9.0005
R6630 iovss.n1617 iovss.n1583 9.0005
R6631 iovss.n1617 iovss.n1560 9.0005
R6632 iovss.n1617 iovss.n1585 9.0005
R6633 iovss.n1617 iovss.n1559 9.0005
R6634 iovss.n1617 iovss.n1587 9.0005
R6635 iovss.n1617 iovss.n1558 9.0005
R6636 iovss.n1617 iovss.n1589 9.0005
R6637 iovss.n1617 iovss.n1557 9.0005
R6638 iovss.n1617 iovss.n1591 9.0005
R6639 iovss.n1617 iovss.n1556 9.0005
R6640 iovss.n1617 iovss.n1593 9.0005
R6641 iovss.n1617 iovss.n1555 9.0005
R6642 iovss.n1617 iovss.n1595 9.0005
R6643 iovss.n1617 iovss.n1554 9.0005
R6644 iovss.n1617 iovss.n1596 9.0005
R6645 iovss.n1617 iovss.n1553 9.0005
R6646 iovss.n1617 iovss.n1598 9.0005
R6647 iovss.n1617 iovss.n1552 9.0005
R6648 iovss.n1617 iovss.n1599 9.0005
R6649 iovss.n1617 iovss.n1551 9.0005
R6650 iovss.n2396 iovss.n1617 9.0005
R6651 iovss.n2394 iovss.n1617 9.0005
R6652 iovss.n1634 iovss.n1569 9.0005
R6653 iovss.n1634 iovss.n1567 9.0005
R6654 iovss.n1634 iovss.n1571 9.0005
R6655 iovss.n1634 iovss.n1566 9.0005
R6656 iovss.n1634 iovss.n1573 9.0005
R6657 iovss.n1634 iovss.n1565 9.0005
R6658 iovss.n1634 iovss.n1575 9.0005
R6659 iovss.n1634 iovss.n1564 9.0005
R6660 iovss.n1634 iovss.n1577 9.0005
R6661 iovss.n1634 iovss.n1563 9.0005
R6662 iovss.n1634 iovss.n1579 9.0005
R6663 iovss.n1634 iovss.n1562 9.0005
R6664 iovss.n1634 iovss.n1581 9.0005
R6665 iovss.n1634 iovss.n1561 9.0005
R6666 iovss.n1634 iovss.n1583 9.0005
R6667 iovss.n1634 iovss.n1560 9.0005
R6668 iovss.n1634 iovss.n1585 9.0005
R6669 iovss.n1634 iovss.n1559 9.0005
R6670 iovss.n1634 iovss.n1587 9.0005
R6671 iovss.n1634 iovss.n1558 9.0005
R6672 iovss.n1634 iovss.n1589 9.0005
R6673 iovss.n1634 iovss.n1557 9.0005
R6674 iovss.n1634 iovss.n1591 9.0005
R6675 iovss.n1634 iovss.n1556 9.0005
R6676 iovss.n1634 iovss.n1593 9.0005
R6677 iovss.n1634 iovss.n1555 9.0005
R6678 iovss.n1634 iovss.n1595 9.0005
R6679 iovss.n1634 iovss.n1554 9.0005
R6680 iovss.n1634 iovss.n1596 9.0005
R6681 iovss.n1634 iovss.n1553 9.0005
R6682 iovss.n1634 iovss.n1598 9.0005
R6683 iovss.n1634 iovss.n1552 9.0005
R6684 iovss.n1634 iovss.n1599 9.0005
R6685 iovss.n1634 iovss.n1551 9.0005
R6686 iovss.n2396 iovss.n1634 9.0005
R6687 iovss.n2394 iovss.n1634 9.0005
R6688 iovss.n1616 iovss.n1569 9.0005
R6689 iovss.n1616 iovss.n1567 9.0005
R6690 iovss.n1616 iovss.n1571 9.0005
R6691 iovss.n1616 iovss.n1566 9.0005
R6692 iovss.n1616 iovss.n1573 9.0005
R6693 iovss.n1616 iovss.n1565 9.0005
R6694 iovss.n1616 iovss.n1575 9.0005
R6695 iovss.n1616 iovss.n1564 9.0005
R6696 iovss.n1616 iovss.n1577 9.0005
R6697 iovss.n1616 iovss.n1563 9.0005
R6698 iovss.n1616 iovss.n1579 9.0005
R6699 iovss.n1616 iovss.n1562 9.0005
R6700 iovss.n1616 iovss.n1581 9.0005
R6701 iovss.n1616 iovss.n1561 9.0005
R6702 iovss.n1616 iovss.n1583 9.0005
R6703 iovss.n1616 iovss.n1560 9.0005
R6704 iovss.n1616 iovss.n1585 9.0005
R6705 iovss.n1616 iovss.n1559 9.0005
R6706 iovss.n1616 iovss.n1587 9.0005
R6707 iovss.n1616 iovss.n1558 9.0005
R6708 iovss.n1616 iovss.n1589 9.0005
R6709 iovss.n1616 iovss.n1557 9.0005
R6710 iovss.n1616 iovss.n1591 9.0005
R6711 iovss.n1616 iovss.n1556 9.0005
R6712 iovss.n1616 iovss.n1593 9.0005
R6713 iovss.n1616 iovss.n1555 9.0005
R6714 iovss.n1616 iovss.n1595 9.0005
R6715 iovss.n1616 iovss.n1554 9.0005
R6716 iovss.n1616 iovss.n1596 9.0005
R6717 iovss.n1616 iovss.n1553 9.0005
R6718 iovss.n1616 iovss.n1598 9.0005
R6719 iovss.n1616 iovss.n1552 9.0005
R6720 iovss.n1616 iovss.n1599 9.0005
R6721 iovss.n1616 iovss.n1551 9.0005
R6722 iovss.n2396 iovss.n1616 9.0005
R6723 iovss.n2394 iovss.n1616 9.0005
R6724 iovss.n1635 iovss.n1569 9.0005
R6725 iovss.n1635 iovss.n1567 9.0005
R6726 iovss.n1635 iovss.n1571 9.0005
R6727 iovss.n1635 iovss.n1566 9.0005
R6728 iovss.n1635 iovss.n1573 9.0005
R6729 iovss.n1635 iovss.n1565 9.0005
R6730 iovss.n1635 iovss.n1575 9.0005
R6731 iovss.n1635 iovss.n1564 9.0005
R6732 iovss.n1635 iovss.n1577 9.0005
R6733 iovss.n1635 iovss.n1563 9.0005
R6734 iovss.n1635 iovss.n1579 9.0005
R6735 iovss.n1635 iovss.n1562 9.0005
R6736 iovss.n1635 iovss.n1581 9.0005
R6737 iovss.n1635 iovss.n1561 9.0005
R6738 iovss.n1635 iovss.n1583 9.0005
R6739 iovss.n1635 iovss.n1560 9.0005
R6740 iovss.n1635 iovss.n1585 9.0005
R6741 iovss.n1635 iovss.n1559 9.0005
R6742 iovss.n1635 iovss.n1587 9.0005
R6743 iovss.n1635 iovss.n1558 9.0005
R6744 iovss.n1635 iovss.n1589 9.0005
R6745 iovss.n1635 iovss.n1557 9.0005
R6746 iovss.n1635 iovss.n1591 9.0005
R6747 iovss.n1635 iovss.n1556 9.0005
R6748 iovss.n1635 iovss.n1593 9.0005
R6749 iovss.n1635 iovss.n1555 9.0005
R6750 iovss.n1635 iovss.n1595 9.0005
R6751 iovss.n1635 iovss.n1554 9.0005
R6752 iovss.n1635 iovss.n1596 9.0005
R6753 iovss.n1635 iovss.n1553 9.0005
R6754 iovss.n1635 iovss.n1598 9.0005
R6755 iovss.n1635 iovss.n1552 9.0005
R6756 iovss.n1635 iovss.n1599 9.0005
R6757 iovss.n1635 iovss.n1551 9.0005
R6758 iovss.n2396 iovss.n1635 9.0005
R6759 iovss.n2394 iovss.n1635 9.0005
R6760 iovss.n1615 iovss.n1569 9.0005
R6761 iovss.n1615 iovss.n1567 9.0005
R6762 iovss.n1615 iovss.n1571 9.0005
R6763 iovss.n1615 iovss.n1566 9.0005
R6764 iovss.n1615 iovss.n1573 9.0005
R6765 iovss.n1615 iovss.n1565 9.0005
R6766 iovss.n1615 iovss.n1575 9.0005
R6767 iovss.n1615 iovss.n1564 9.0005
R6768 iovss.n1615 iovss.n1577 9.0005
R6769 iovss.n1615 iovss.n1563 9.0005
R6770 iovss.n1615 iovss.n1579 9.0005
R6771 iovss.n1615 iovss.n1562 9.0005
R6772 iovss.n1615 iovss.n1581 9.0005
R6773 iovss.n1615 iovss.n1561 9.0005
R6774 iovss.n1615 iovss.n1583 9.0005
R6775 iovss.n1615 iovss.n1560 9.0005
R6776 iovss.n1615 iovss.n1585 9.0005
R6777 iovss.n1615 iovss.n1559 9.0005
R6778 iovss.n1615 iovss.n1587 9.0005
R6779 iovss.n1615 iovss.n1558 9.0005
R6780 iovss.n1615 iovss.n1589 9.0005
R6781 iovss.n1615 iovss.n1557 9.0005
R6782 iovss.n1615 iovss.n1591 9.0005
R6783 iovss.n1615 iovss.n1556 9.0005
R6784 iovss.n1615 iovss.n1593 9.0005
R6785 iovss.n1615 iovss.n1555 9.0005
R6786 iovss.n1615 iovss.n1595 9.0005
R6787 iovss.n1615 iovss.n1554 9.0005
R6788 iovss.n1615 iovss.n1596 9.0005
R6789 iovss.n1615 iovss.n1553 9.0005
R6790 iovss.n1615 iovss.n1598 9.0005
R6791 iovss.n1615 iovss.n1552 9.0005
R6792 iovss.n1615 iovss.n1599 9.0005
R6793 iovss.n1615 iovss.n1551 9.0005
R6794 iovss.n2396 iovss.n1615 9.0005
R6795 iovss.n2394 iovss.n1615 9.0005
R6796 iovss.n1636 iovss.n1569 9.0005
R6797 iovss.n1636 iovss.n1567 9.0005
R6798 iovss.n1636 iovss.n1571 9.0005
R6799 iovss.n1636 iovss.n1566 9.0005
R6800 iovss.n1636 iovss.n1573 9.0005
R6801 iovss.n1636 iovss.n1565 9.0005
R6802 iovss.n1636 iovss.n1575 9.0005
R6803 iovss.n1636 iovss.n1564 9.0005
R6804 iovss.n1636 iovss.n1577 9.0005
R6805 iovss.n1636 iovss.n1563 9.0005
R6806 iovss.n1636 iovss.n1579 9.0005
R6807 iovss.n1636 iovss.n1562 9.0005
R6808 iovss.n1636 iovss.n1581 9.0005
R6809 iovss.n1636 iovss.n1561 9.0005
R6810 iovss.n1636 iovss.n1583 9.0005
R6811 iovss.n1636 iovss.n1560 9.0005
R6812 iovss.n1636 iovss.n1585 9.0005
R6813 iovss.n1636 iovss.n1559 9.0005
R6814 iovss.n1636 iovss.n1587 9.0005
R6815 iovss.n1636 iovss.n1558 9.0005
R6816 iovss.n1636 iovss.n1589 9.0005
R6817 iovss.n1636 iovss.n1557 9.0005
R6818 iovss.n1636 iovss.n1591 9.0005
R6819 iovss.n1636 iovss.n1556 9.0005
R6820 iovss.n1636 iovss.n1593 9.0005
R6821 iovss.n1636 iovss.n1555 9.0005
R6822 iovss.n1636 iovss.n1595 9.0005
R6823 iovss.n1636 iovss.n1554 9.0005
R6824 iovss.n1636 iovss.n1596 9.0005
R6825 iovss.n1636 iovss.n1553 9.0005
R6826 iovss.n1636 iovss.n1598 9.0005
R6827 iovss.n1636 iovss.n1552 9.0005
R6828 iovss.n1636 iovss.n1599 9.0005
R6829 iovss.n1636 iovss.n1551 9.0005
R6830 iovss.n2396 iovss.n1636 9.0005
R6831 iovss.n2394 iovss.n1636 9.0005
R6832 iovss.n1614 iovss.n1569 9.0005
R6833 iovss.n1614 iovss.n1567 9.0005
R6834 iovss.n1614 iovss.n1571 9.0005
R6835 iovss.n1614 iovss.n1566 9.0005
R6836 iovss.n1614 iovss.n1573 9.0005
R6837 iovss.n1614 iovss.n1565 9.0005
R6838 iovss.n1614 iovss.n1575 9.0005
R6839 iovss.n1614 iovss.n1564 9.0005
R6840 iovss.n1614 iovss.n1577 9.0005
R6841 iovss.n1614 iovss.n1563 9.0005
R6842 iovss.n1614 iovss.n1579 9.0005
R6843 iovss.n1614 iovss.n1562 9.0005
R6844 iovss.n1614 iovss.n1581 9.0005
R6845 iovss.n1614 iovss.n1561 9.0005
R6846 iovss.n1614 iovss.n1583 9.0005
R6847 iovss.n1614 iovss.n1560 9.0005
R6848 iovss.n1614 iovss.n1585 9.0005
R6849 iovss.n1614 iovss.n1559 9.0005
R6850 iovss.n1614 iovss.n1587 9.0005
R6851 iovss.n1614 iovss.n1558 9.0005
R6852 iovss.n1614 iovss.n1589 9.0005
R6853 iovss.n1614 iovss.n1557 9.0005
R6854 iovss.n1614 iovss.n1591 9.0005
R6855 iovss.n1614 iovss.n1556 9.0005
R6856 iovss.n1614 iovss.n1593 9.0005
R6857 iovss.n1614 iovss.n1555 9.0005
R6858 iovss.n1614 iovss.n1595 9.0005
R6859 iovss.n1614 iovss.n1554 9.0005
R6860 iovss.n1614 iovss.n1596 9.0005
R6861 iovss.n1614 iovss.n1553 9.0005
R6862 iovss.n1614 iovss.n1598 9.0005
R6863 iovss.n1614 iovss.n1552 9.0005
R6864 iovss.n1614 iovss.n1599 9.0005
R6865 iovss.n1614 iovss.n1551 9.0005
R6866 iovss.n2396 iovss.n1614 9.0005
R6867 iovss.n2394 iovss.n1614 9.0005
R6868 iovss.n1637 iovss.n1569 9.0005
R6869 iovss.n1637 iovss.n1567 9.0005
R6870 iovss.n1637 iovss.n1571 9.0005
R6871 iovss.n1637 iovss.n1566 9.0005
R6872 iovss.n1637 iovss.n1573 9.0005
R6873 iovss.n1637 iovss.n1565 9.0005
R6874 iovss.n1637 iovss.n1575 9.0005
R6875 iovss.n1637 iovss.n1564 9.0005
R6876 iovss.n1637 iovss.n1577 9.0005
R6877 iovss.n1637 iovss.n1563 9.0005
R6878 iovss.n1637 iovss.n1579 9.0005
R6879 iovss.n1637 iovss.n1562 9.0005
R6880 iovss.n1637 iovss.n1581 9.0005
R6881 iovss.n1637 iovss.n1561 9.0005
R6882 iovss.n1637 iovss.n1583 9.0005
R6883 iovss.n1637 iovss.n1560 9.0005
R6884 iovss.n1637 iovss.n1585 9.0005
R6885 iovss.n1637 iovss.n1559 9.0005
R6886 iovss.n1637 iovss.n1587 9.0005
R6887 iovss.n1637 iovss.n1558 9.0005
R6888 iovss.n1637 iovss.n1589 9.0005
R6889 iovss.n1637 iovss.n1557 9.0005
R6890 iovss.n1637 iovss.n1591 9.0005
R6891 iovss.n1637 iovss.n1556 9.0005
R6892 iovss.n1637 iovss.n1593 9.0005
R6893 iovss.n1637 iovss.n1555 9.0005
R6894 iovss.n1637 iovss.n1595 9.0005
R6895 iovss.n1637 iovss.n1554 9.0005
R6896 iovss.n1637 iovss.n1596 9.0005
R6897 iovss.n1637 iovss.n1553 9.0005
R6898 iovss.n1637 iovss.n1598 9.0005
R6899 iovss.n1637 iovss.n1552 9.0005
R6900 iovss.n1637 iovss.n1599 9.0005
R6901 iovss.n1637 iovss.n1551 9.0005
R6902 iovss.n2396 iovss.n1637 9.0005
R6903 iovss.n2394 iovss.n1637 9.0005
R6904 iovss.n1613 iovss.n1569 9.0005
R6905 iovss.n1613 iovss.n1567 9.0005
R6906 iovss.n1613 iovss.n1571 9.0005
R6907 iovss.n1613 iovss.n1566 9.0005
R6908 iovss.n1613 iovss.n1573 9.0005
R6909 iovss.n1613 iovss.n1565 9.0005
R6910 iovss.n1613 iovss.n1575 9.0005
R6911 iovss.n1613 iovss.n1564 9.0005
R6912 iovss.n1613 iovss.n1577 9.0005
R6913 iovss.n1613 iovss.n1563 9.0005
R6914 iovss.n1613 iovss.n1579 9.0005
R6915 iovss.n1613 iovss.n1562 9.0005
R6916 iovss.n1613 iovss.n1581 9.0005
R6917 iovss.n1613 iovss.n1561 9.0005
R6918 iovss.n1613 iovss.n1583 9.0005
R6919 iovss.n1613 iovss.n1560 9.0005
R6920 iovss.n1613 iovss.n1585 9.0005
R6921 iovss.n1613 iovss.n1559 9.0005
R6922 iovss.n1613 iovss.n1587 9.0005
R6923 iovss.n1613 iovss.n1558 9.0005
R6924 iovss.n1613 iovss.n1589 9.0005
R6925 iovss.n1613 iovss.n1557 9.0005
R6926 iovss.n1613 iovss.n1591 9.0005
R6927 iovss.n1613 iovss.n1556 9.0005
R6928 iovss.n1613 iovss.n1593 9.0005
R6929 iovss.n1613 iovss.n1555 9.0005
R6930 iovss.n1613 iovss.n1595 9.0005
R6931 iovss.n1613 iovss.n1554 9.0005
R6932 iovss.n1613 iovss.n1596 9.0005
R6933 iovss.n1613 iovss.n1553 9.0005
R6934 iovss.n1613 iovss.n1598 9.0005
R6935 iovss.n1613 iovss.n1552 9.0005
R6936 iovss.n1613 iovss.n1599 9.0005
R6937 iovss.n1613 iovss.n1551 9.0005
R6938 iovss.n2396 iovss.n1613 9.0005
R6939 iovss.n2394 iovss.n1613 9.0005
R6940 iovss.n1638 iovss.n1569 9.0005
R6941 iovss.n1638 iovss.n1567 9.0005
R6942 iovss.n1638 iovss.n1571 9.0005
R6943 iovss.n1638 iovss.n1566 9.0005
R6944 iovss.n1638 iovss.n1573 9.0005
R6945 iovss.n1638 iovss.n1565 9.0005
R6946 iovss.n1638 iovss.n1575 9.0005
R6947 iovss.n1638 iovss.n1564 9.0005
R6948 iovss.n1638 iovss.n1577 9.0005
R6949 iovss.n1638 iovss.n1563 9.0005
R6950 iovss.n1638 iovss.n1579 9.0005
R6951 iovss.n1638 iovss.n1562 9.0005
R6952 iovss.n1638 iovss.n1581 9.0005
R6953 iovss.n1638 iovss.n1561 9.0005
R6954 iovss.n1638 iovss.n1583 9.0005
R6955 iovss.n1638 iovss.n1560 9.0005
R6956 iovss.n1638 iovss.n1585 9.0005
R6957 iovss.n1638 iovss.n1559 9.0005
R6958 iovss.n1638 iovss.n1587 9.0005
R6959 iovss.n1638 iovss.n1558 9.0005
R6960 iovss.n1638 iovss.n1589 9.0005
R6961 iovss.n1638 iovss.n1557 9.0005
R6962 iovss.n1638 iovss.n1591 9.0005
R6963 iovss.n1638 iovss.n1556 9.0005
R6964 iovss.n1638 iovss.n1593 9.0005
R6965 iovss.n1638 iovss.n1555 9.0005
R6966 iovss.n1638 iovss.n1595 9.0005
R6967 iovss.n1638 iovss.n1554 9.0005
R6968 iovss.n1638 iovss.n1596 9.0005
R6969 iovss.n1638 iovss.n1553 9.0005
R6970 iovss.n1638 iovss.n1598 9.0005
R6971 iovss.n1638 iovss.n1552 9.0005
R6972 iovss.n1638 iovss.n1599 9.0005
R6973 iovss.n1638 iovss.n1551 9.0005
R6974 iovss.n2396 iovss.n1638 9.0005
R6975 iovss.n2394 iovss.n1638 9.0005
R6976 iovss.n1612 iovss.n1569 9.0005
R6977 iovss.n1612 iovss.n1567 9.0005
R6978 iovss.n1612 iovss.n1571 9.0005
R6979 iovss.n1612 iovss.n1566 9.0005
R6980 iovss.n1612 iovss.n1573 9.0005
R6981 iovss.n1612 iovss.n1565 9.0005
R6982 iovss.n1612 iovss.n1575 9.0005
R6983 iovss.n1612 iovss.n1564 9.0005
R6984 iovss.n1612 iovss.n1577 9.0005
R6985 iovss.n1612 iovss.n1563 9.0005
R6986 iovss.n1612 iovss.n1579 9.0005
R6987 iovss.n1612 iovss.n1562 9.0005
R6988 iovss.n1612 iovss.n1581 9.0005
R6989 iovss.n1612 iovss.n1561 9.0005
R6990 iovss.n1612 iovss.n1583 9.0005
R6991 iovss.n1612 iovss.n1560 9.0005
R6992 iovss.n1612 iovss.n1585 9.0005
R6993 iovss.n1612 iovss.n1559 9.0005
R6994 iovss.n1612 iovss.n1587 9.0005
R6995 iovss.n1612 iovss.n1558 9.0005
R6996 iovss.n1612 iovss.n1589 9.0005
R6997 iovss.n1612 iovss.n1557 9.0005
R6998 iovss.n1612 iovss.n1591 9.0005
R6999 iovss.n1612 iovss.n1556 9.0005
R7000 iovss.n1612 iovss.n1593 9.0005
R7001 iovss.n1612 iovss.n1555 9.0005
R7002 iovss.n1612 iovss.n1595 9.0005
R7003 iovss.n1612 iovss.n1554 9.0005
R7004 iovss.n1612 iovss.n1596 9.0005
R7005 iovss.n1612 iovss.n1553 9.0005
R7006 iovss.n1612 iovss.n1598 9.0005
R7007 iovss.n1612 iovss.n1552 9.0005
R7008 iovss.n1612 iovss.n1599 9.0005
R7009 iovss.n1612 iovss.n1551 9.0005
R7010 iovss.n2396 iovss.n1612 9.0005
R7011 iovss.n2394 iovss.n1612 9.0005
R7012 iovss.n1639 iovss.n1569 9.0005
R7013 iovss.n1639 iovss.n1567 9.0005
R7014 iovss.n1639 iovss.n1571 9.0005
R7015 iovss.n1639 iovss.n1566 9.0005
R7016 iovss.n1639 iovss.n1573 9.0005
R7017 iovss.n1639 iovss.n1565 9.0005
R7018 iovss.n1639 iovss.n1575 9.0005
R7019 iovss.n1639 iovss.n1564 9.0005
R7020 iovss.n1639 iovss.n1577 9.0005
R7021 iovss.n1639 iovss.n1563 9.0005
R7022 iovss.n1639 iovss.n1579 9.0005
R7023 iovss.n1639 iovss.n1562 9.0005
R7024 iovss.n1639 iovss.n1581 9.0005
R7025 iovss.n1639 iovss.n1561 9.0005
R7026 iovss.n1639 iovss.n1583 9.0005
R7027 iovss.n1639 iovss.n1560 9.0005
R7028 iovss.n1639 iovss.n1585 9.0005
R7029 iovss.n1639 iovss.n1559 9.0005
R7030 iovss.n1639 iovss.n1587 9.0005
R7031 iovss.n1639 iovss.n1558 9.0005
R7032 iovss.n1639 iovss.n1589 9.0005
R7033 iovss.n1639 iovss.n1557 9.0005
R7034 iovss.n1639 iovss.n1591 9.0005
R7035 iovss.n1639 iovss.n1556 9.0005
R7036 iovss.n1639 iovss.n1593 9.0005
R7037 iovss.n1639 iovss.n1555 9.0005
R7038 iovss.n1639 iovss.n1595 9.0005
R7039 iovss.n1639 iovss.n1554 9.0005
R7040 iovss.n1639 iovss.n1596 9.0005
R7041 iovss.n1639 iovss.n1553 9.0005
R7042 iovss.n1639 iovss.n1598 9.0005
R7043 iovss.n1639 iovss.n1552 9.0005
R7044 iovss.n1639 iovss.n1599 9.0005
R7045 iovss.n1639 iovss.n1551 9.0005
R7046 iovss.n2396 iovss.n1639 9.0005
R7047 iovss.n2394 iovss.n1639 9.0005
R7048 iovss.n1611 iovss.n1569 9.0005
R7049 iovss.n1611 iovss.n1567 9.0005
R7050 iovss.n1611 iovss.n1571 9.0005
R7051 iovss.n1611 iovss.n1566 9.0005
R7052 iovss.n1611 iovss.n1573 9.0005
R7053 iovss.n1611 iovss.n1565 9.0005
R7054 iovss.n1611 iovss.n1575 9.0005
R7055 iovss.n1611 iovss.n1564 9.0005
R7056 iovss.n1611 iovss.n1577 9.0005
R7057 iovss.n1611 iovss.n1563 9.0005
R7058 iovss.n1611 iovss.n1579 9.0005
R7059 iovss.n1611 iovss.n1562 9.0005
R7060 iovss.n1611 iovss.n1581 9.0005
R7061 iovss.n1611 iovss.n1561 9.0005
R7062 iovss.n1611 iovss.n1583 9.0005
R7063 iovss.n1611 iovss.n1560 9.0005
R7064 iovss.n1611 iovss.n1585 9.0005
R7065 iovss.n1611 iovss.n1559 9.0005
R7066 iovss.n1611 iovss.n1587 9.0005
R7067 iovss.n1611 iovss.n1558 9.0005
R7068 iovss.n1611 iovss.n1589 9.0005
R7069 iovss.n1611 iovss.n1557 9.0005
R7070 iovss.n1611 iovss.n1591 9.0005
R7071 iovss.n1611 iovss.n1556 9.0005
R7072 iovss.n1611 iovss.n1593 9.0005
R7073 iovss.n1611 iovss.n1555 9.0005
R7074 iovss.n1611 iovss.n1595 9.0005
R7075 iovss.n1611 iovss.n1554 9.0005
R7076 iovss.n1611 iovss.n1596 9.0005
R7077 iovss.n1611 iovss.n1553 9.0005
R7078 iovss.n1611 iovss.n1598 9.0005
R7079 iovss.n1611 iovss.n1552 9.0005
R7080 iovss.n1611 iovss.n1599 9.0005
R7081 iovss.n1611 iovss.n1551 9.0005
R7082 iovss.n2396 iovss.n1611 9.0005
R7083 iovss.n2394 iovss.n1611 9.0005
R7084 iovss.n1640 iovss.n1569 9.0005
R7085 iovss.n1640 iovss.n1567 9.0005
R7086 iovss.n1640 iovss.n1571 9.0005
R7087 iovss.n1640 iovss.n1566 9.0005
R7088 iovss.n1640 iovss.n1573 9.0005
R7089 iovss.n1640 iovss.n1565 9.0005
R7090 iovss.n1640 iovss.n1575 9.0005
R7091 iovss.n1640 iovss.n1564 9.0005
R7092 iovss.n1640 iovss.n1577 9.0005
R7093 iovss.n1640 iovss.n1563 9.0005
R7094 iovss.n1640 iovss.n1579 9.0005
R7095 iovss.n1640 iovss.n1562 9.0005
R7096 iovss.n1640 iovss.n1581 9.0005
R7097 iovss.n1640 iovss.n1561 9.0005
R7098 iovss.n1640 iovss.n1583 9.0005
R7099 iovss.n1640 iovss.n1560 9.0005
R7100 iovss.n1640 iovss.n1585 9.0005
R7101 iovss.n1640 iovss.n1559 9.0005
R7102 iovss.n1640 iovss.n1587 9.0005
R7103 iovss.n1640 iovss.n1558 9.0005
R7104 iovss.n1640 iovss.n1589 9.0005
R7105 iovss.n1640 iovss.n1557 9.0005
R7106 iovss.n1640 iovss.n1591 9.0005
R7107 iovss.n1640 iovss.n1556 9.0005
R7108 iovss.n1640 iovss.n1593 9.0005
R7109 iovss.n1640 iovss.n1555 9.0005
R7110 iovss.n1640 iovss.n1595 9.0005
R7111 iovss.n1640 iovss.n1554 9.0005
R7112 iovss.n1640 iovss.n1596 9.0005
R7113 iovss.n1640 iovss.n1553 9.0005
R7114 iovss.n1640 iovss.n1598 9.0005
R7115 iovss.n1640 iovss.n1552 9.0005
R7116 iovss.n1640 iovss.n1599 9.0005
R7117 iovss.n1640 iovss.n1551 9.0005
R7118 iovss.n2396 iovss.n1640 9.0005
R7119 iovss.n2394 iovss.n1640 9.0005
R7120 iovss.n1610 iovss.n1569 9.0005
R7121 iovss.n1610 iovss.n1567 9.0005
R7122 iovss.n1610 iovss.n1571 9.0005
R7123 iovss.n1610 iovss.n1566 9.0005
R7124 iovss.n1610 iovss.n1573 9.0005
R7125 iovss.n1610 iovss.n1565 9.0005
R7126 iovss.n1610 iovss.n1575 9.0005
R7127 iovss.n1610 iovss.n1564 9.0005
R7128 iovss.n1610 iovss.n1577 9.0005
R7129 iovss.n1610 iovss.n1563 9.0005
R7130 iovss.n1610 iovss.n1579 9.0005
R7131 iovss.n1610 iovss.n1562 9.0005
R7132 iovss.n1610 iovss.n1581 9.0005
R7133 iovss.n1610 iovss.n1561 9.0005
R7134 iovss.n1610 iovss.n1583 9.0005
R7135 iovss.n1610 iovss.n1560 9.0005
R7136 iovss.n1610 iovss.n1585 9.0005
R7137 iovss.n1610 iovss.n1559 9.0005
R7138 iovss.n1610 iovss.n1587 9.0005
R7139 iovss.n1610 iovss.n1558 9.0005
R7140 iovss.n1610 iovss.n1589 9.0005
R7141 iovss.n1610 iovss.n1557 9.0005
R7142 iovss.n1610 iovss.n1591 9.0005
R7143 iovss.n1610 iovss.n1556 9.0005
R7144 iovss.n1610 iovss.n1593 9.0005
R7145 iovss.n1610 iovss.n1555 9.0005
R7146 iovss.n1610 iovss.n1595 9.0005
R7147 iovss.n1610 iovss.n1554 9.0005
R7148 iovss.n1610 iovss.n1596 9.0005
R7149 iovss.n1610 iovss.n1553 9.0005
R7150 iovss.n1610 iovss.n1598 9.0005
R7151 iovss.n1610 iovss.n1552 9.0005
R7152 iovss.n1610 iovss.n1599 9.0005
R7153 iovss.n1610 iovss.n1551 9.0005
R7154 iovss.n2396 iovss.n1610 9.0005
R7155 iovss.n2394 iovss.n1610 9.0005
R7156 iovss.n1641 iovss.n1569 9.0005
R7157 iovss.n1641 iovss.n1567 9.0005
R7158 iovss.n1641 iovss.n1571 9.0005
R7159 iovss.n1641 iovss.n1566 9.0005
R7160 iovss.n1641 iovss.n1573 9.0005
R7161 iovss.n1641 iovss.n1565 9.0005
R7162 iovss.n1641 iovss.n1575 9.0005
R7163 iovss.n1641 iovss.n1564 9.0005
R7164 iovss.n1641 iovss.n1577 9.0005
R7165 iovss.n1641 iovss.n1563 9.0005
R7166 iovss.n1641 iovss.n1579 9.0005
R7167 iovss.n1641 iovss.n1562 9.0005
R7168 iovss.n1641 iovss.n1581 9.0005
R7169 iovss.n1641 iovss.n1561 9.0005
R7170 iovss.n1641 iovss.n1583 9.0005
R7171 iovss.n1641 iovss.n1560 9.0005
R7172 iovss.n1641 iovss.n1585 9.0005
R7173 iovss.n1641 iovss.n1559 9.0005
R7174 iovss.n1641 iovss.n1587 9.0005
R7175 iovss.n1641 iovss.n1558 9.0005
R7176 iovss.n1641 iovss.n1589 9.0005
R7177 iovss.n1641 iovss.n1557 9.0005
R7178 iovss.n1641 iovss.n1591 9.0005
R7179 iovss.n1641 iovss.n1556 9.0005
R7180 iovss.n1641 iovss.n1593 9.0005
R7181 iovss.n1641 iovss.n1555 9.0005
R7182 iovss.n1641 iovss.n1595 9.0005
R7183 iovss.n1641 iovss.n1554 9.0005
R7184 iovss.n1641 iovss.n1596 9.0005
R7185 iovss.n1641 iovss.n1553 9.0005
R7186 iovss.n1641 iovss.n1598 9.0005
R7187 iovss.n1641 iovss.n1552 9.0005
R7188 iovss.n1641 iovss.n1599 9.0005
R7189 iovss.n1641 iovss.n1551 9.0005
R7190 iovss.n2396 iovss.n1641 9.0005
R7191 iovss.n2394 iovss.n1641 9.0005
R7192 iovss.n1609 iovss.n1569 9.0005
R7193 iovss.n1609 iovss.n1567 9.0005
R7194 iovss.n1609 iovss.n1571 9.0005
R7195 iovss.n1609 iovss.n1566 9.0005
R7196 iovss.n1609 iovss.n1573 9.0005
R7197 iovss.n1609 iovss.n1565 9.0005
R7198 iovss.n1609 iovss.n1575 9.0005
R7199 iovss.n1609 iovss.n1564 9.0005
R7200 iovss.n1609 iovss.n1577 9.0005
R7201 iovss.n1609 iovss.n1563 9.0005
R7202 iovss.n1609 iovss.n1579 9.0005
R7203 iovss.n1609 iovss.n1562 9.0005
R7204 iovss.n1609 iovss.n1581 9.0005
R7205 iovss.n1609 iovss.n1561 9.0005
R7206 iovss.n1609 iovss.n1583 9.0005
R7207 iovss.n1609 iovss.n1560 9.0005
R7208 iovss.n1609 iovss.n1585 9.0005
R7209 iovss.n1609 iovss.n1559 9.0005
R7210 iovss.n1609 iovss.n1587 9.0005
R7211 iovss.n1609 iovss.n1558 9.0005
R7212 iovss.n1609 iovss.n1589 9.0005
R7213 iovss.n1609 iovss.n1557 9.0005
R7214 iovss.n1609 iovss.n1591 9.0005
R7215 iovss.n1609 iovss.n1556 9.0005
R7216 iovss.n1609 iovss.n1593 9.0005
R7217 iovss.n1609 iovss.n1555 9.0005
R7218 iovss.n1609 iovss.n1595 9.0005
R7219 iovss.n1609 iovss.n1554 9.0005
R7220 iovss.n1609 iovss.n1596 9.0005
R7221 iovss.n1609 iovss.n1553 9.0005
R7222 iovss.n1609 iovss.n1598 9.0005
R7223 iovss.n1609 iovss.n1552 9.0005
R7224 iovss.n1609 iovss.n1599 9.0005
R7225 iovss.n1609 iovss.n1551 9.0005
R7226 iovss.n2396 iovss.n1609 9.0005
R7227 iovss.n2394 iovss.n1609 9.0005
R7228 iovss.n1642 iovss.n1569 9.0005
R7229 iovss.n1642 iovss.n1567 9.0005
R7230 iovss.n1642 iovss.n1571 9.0005
R7231 iovss.n1642 iovss.n1566 9.0005
R7232 iovss.n1642 iovss.n1573 9.0005
R7233 iovss.n1642 iovss.n1565 9.0005
R7234 iovss.n1642 iovss.n1575 9.0005
R7235 iovss.n1642 iovss.n1564 9.0005
R7236 iovss.n1642 iovss.n1577 9.0005
R7237 iovss.n1642 iovss.n1563 9.0005
R7238 iovss.n1642 iovss.n1579 9.0005
R7239 iovss.n1642 iovss.n1562 9.0005
R7240 iovss.n1642 iovss.n1581 9.0005
R7241 iovss.n1642 iovss.n1561 9.0005
R7242 iovss.n1642 iovss.n1583 9.0005
R7243 iovss.n1642 iovss.n1560 9.0005
R7244 iovss.n1642 iovss.n1585 9.0005
R7245 iovss.n1642 iovss.n1559 9.0005
R7246 iovss.n1642 iovss.n1587 9.0005
R7247 iovss.n1642 iovss.n1558 9.0005
R7248 iovss.n1642 iovss.n1589 9.0005
R7249 iovss.n1642 iovss.n1557 9.0005
R7250 iovss.n1642 iovss.n1591 9.0005
R7251 iovss.n1642 iovss.n1556 9.0005
R7252 iovss.n1642 iovss.n1593 9.0005
R7253 iovss.n1642 iovss.n1555 9.0005
R7254 iovss.n1642 iovss.n1595 9.0005
R7255 iovss.n1642 iovss.n1554 9.0005
R7256 iovss.n1642 iovss.n1596 9.0005
R7257 iovss.n1642 iovss.n1553 9.0005
R7258 iovss.n1642 iovss.n1598 9.0005
R7259 iovss.n1642 iovss.n1552 9.0005
R7260 iovss.n1642 iovss.n1599 9.0005
R7261 iovss.n1642 iovss.n1551 9.0005
R7262 iovss.n2396 iovss.n1642 9.0005
R7263 iovss.n2394 iovss.n1642 9.0005
R7264 iovss.n1608 iovss.n1569 9.0005
R7265 iovss.n1608 iovss.n1567 9.0005
R7266 iovss.n1608 iovss.n1571 9.0005
R7267 iovss.n1608 iovss.n1566 9.0005
R7268 iovss.n1608 iovss.n1573 9.0005
R7269 iovss.n1608 iovss.n1565 9.0005
R7270 iovss.n1608 iovss.n1575 9.0005
R7271 iovss.n1608 iovss.n1564 9.0005
R7272 iovss.n1608 iovss.n1577 9.0005
R7273 iovss.n1608 iovss.n1563 9.0005
R7274 iovss.n1608 iovss.n1579 9.0005
R7275 iovss.n1608 iovss.n1562 9.0005
R7276 iovss.n1608 iovss.n1581 9.0005
R7277 iovss.n1608 iovss.n1561 9.0005
R7278 iovss.n1608 iovss.n1583 9.0005
R7279 iovss.n1608 iovss.n1560 9.0005
R7280 iovss.n1608 iovss.n1585 9.0005
R7281 iovss.n1608 iovss.n1559 9.0005
R7282 iovss.n1608 iovss.n1587 9.0005
R7283 iovss.n1608 iovss.n1558 9.0005
R7284 iovss.n1608 iovss.n1589 9.0005
R7285 iovss.n1608 iovss.n1557 9.0005
R7286 iovss.n1608 iovss.n1591 9.0005
R7287 iovss.n1608 iovss.n1556 9.0005
R7288 iovss.n1608 iovss.n1593 9.0005
R7289 iovss.n1608 iovss.n1555 9.0005
R7290 iovss.n1608 iovss.n1595 9.0005
R7291 iovss.n1608 iovss.n1554 9.0005
R7292 iovss.n1608 iovss.n1596 9.0005
R7293 iovss.n1608 iovss.n1553 9.0005
R7294 iovss.n1608 iovss.n1598 9.0005
R7295 iovss.n1608 iovss.n1552 9.0005
R7296 iovss.n1608 iovss.n1599 9.0005
R7297 iovss.n1608 iovss.n1551 9.0005
R7298 iovss.n2396 iovss.n1608 9.0005
R7299 iovss.n2394 iovss.n1608 9.0005
R7300 iovss.n1643 iovss.n1569 9.0005
R7301 iovss.n1643 iovss.n1567 9.0005
R7302 iovss.n1643 iovss.n1571 9.0005
R7303 iovss.n1643 iovss.n1566 9.0005
R7304 iovss.n1643 iovss.n1573 9.0005
R7305 iovss.n1643 iovss.n1565 9.0005
R7306 iovss.n1643 iovss.n1575 9.0005
R7307 iovss.n1643 iovss.n1564 9.0005
R7308 iovss.n1643 iovss.n1577 9.0005
R7309 iovss.n1643 iovss.n1563 9.0005
R7310 iovss.n1643 iovss.n1579 9.0005
R7311 iovss.n1643 iovss.n1562 9.0005
R7312 iovss.n1643 iovss.n1581 9.0005
R7313 iovss.n1643 iovss.n1561 9.0005
R7314 iovss.n1643 iovss.n1583 9.0005
R7315 iovss.n1643 iovss.n1560 9.0005
R7316 iovss.n1643 iovss.n1585 9.0005
R7317 iovss.n1643 iovss.n1559 9.0005
R7318 iovss.n1643 iovss.n1587 9.0005
R7319 iovss.n1643 iovss.n1558 9.0005
R7320 iovss.n1643 iovss.n1589 9.0005
R7321 iovss.n1643 iovss.n1557 9.0005
R7322 iovss.n1643 iovss.n1591 9.0005
R7323 iovss.n1643 iovss.n1556 9.0005
R7324 iovss.n1643 iovss.n1593 9.0005
R7325 iovss.n1643 iovss.n1555 9.0005
R7326 iovss.n1643 iovss.n1595 9.0005
R7327 iovss.n1643 iovss.n1554 9.0005
R7328 iovss.n1643 iovss.n1596 9.0005
R7329 iovss.n1643 iovss.n1553 9.0005
R7330 iovss.n1643 iovss.n1598 9.0005
R7331 iovss.n1643 iovss.n1552 9.0005
R7332 iovss.n1643 iovss.n1599 9.0005
R7333 iovss.n1643 iovss.n1551 9.0005
R7334 iovss.n2396 iovss.n1643 9.0005
R7335 iovss.n2394 iovss.n1643 9.0005
R7336 iovss.n1607 iovss.n1569 9.0005
R7337 iovss.n1607 iovss.n1567 9.0005
R7338 iovss.n1607 iovss.n1571 9.0005
R7339 iovss.n1607 iovss.n1566 9.0005
R7340 iovss.n1607 iovss.n1573 9.0005
R7341 iovss.n1607 iovss.n1565 9.0005
R7342 iovss.n1607 iovss.n1575 9.0005
R7343 iovss.n1607 iovss.n1564 9.0005
R7344 iovss.n1607 iovss.n1577 9.0005
R7345 iovss.n1607 iovss.n1563 9.0005
R7346 iovss.n1607 iovss.n1579 9.0005
R7347 iovss.n1607 iovss.n1562 9.0005
R7348 iovss.n1607 iovss.n1581 9.0005
R7349 iovss.n1607 iovss.n1561 9.0005
R7350 iovss.n1607 iovss.n1583 9.0005
R7351 iovss.n1607 iovss.n1560 9.0005
R7352 iovss.n1607 iovss.n1585 9.0005
R7353 iovss.n1607 iovss.n1559 9.0005
R7354 iovss.n1607 iovss.n1587 9.0005
R7355 iovss.n1607 iovss.n1558 9.0005
R7356 iovss.n1607 iovss.n1589 9.0005
R7357 iovss.n1607 iovss.n1557 9.0005
R7358 iovss.n1607 iovss.n1591 9.0005
R7359 iovss.n1607 iovss.n1556 9.0005
R7360 iovss.n1607 iovss.n1593 9.0005
R7361 iovss.n1607 iovss.n1555 9.0005
R7362 iovss.n1607 iovss.n1595 9.0005
R7363 iovss.n1607 iovss.n1554 9.0005
R7364 iovss.n1607 iovss.n1596 9.0005
R7365 iovss.n1607 iovss.n1553 9.0005
R7366 iovss.n1607 iovss.n1598 9.0005
R7367 iovss.n1607 iovss.n1552 9.0005
R7368 iovss.n1607 iovss.n1599 9.0005
R7369 iovss.n1607 iovss.n1551 9.0005
R7370 iovss.n2396 iovss.n1607 9.0005
R7371 iovss.n2394 iovss.n1607 9.0005
R7372 iovss.n1644 iovss.n1569 9.0005
R7373 iovss.n1644 iovss.n1567 9.0005
R7374 iovss.n1644 iovss.n1571 9.0005
R7375 iovss.n1644 iovss.n1566 9.0005
R7376 iovss.n1644 iovss.n1573 9.0005
R7377 iovss.n1644 iovss.n1565 9.0005
R7378 iovss.n1644 iovss.n1575 9.0005
R7379 iovss.n1644 iovss.n1564 9.0005
R7380 iovss.n1644 iovss.n1577 9.0005
R7381 iovss.n1644 iovss.n1563 9.0005
R7382 iovss.n1644 iovss.n1579 9.0005
R7383 iovss.n1644 iovss.n1562 9.0005
R7384 iovss.n1644 iovss.n1581 9.0005
R7385 iovss.n1644 iovss.n1561 9.0005
R7386 iovss.n1644 iovss.n1583 9.0005
R7387 iovss.n1644 iovss.n1560 9.0005
R7388 iovss.n1644 iovss.n1585 9.0005
R7389 iovss.n1644 iovss.n1559 9.0005
R7390 iovss.n1644 iovss.n1587 9.0005
R7391 iovss.n1644 iovss.n1558 9.0005
R7392 iovss.n1644 iovss.n1589 9.0005
R7393 iovss.n1644 iovss.n1557 9.0005
R7394 iovss.n1644 iovss.n1591 9.0005
R7395 iovss.n1644 iovss.n1556 9.0005
R7396 iovss.n1644 iovss.n1593 9.0005
R7397 iovss.n1644 iovss.n1555 9.0005
R7398 iovss.n1644 iovss.n1595 9.0005
R7399 iovss.n1644 iovss.n1554 9.0005
R7400 iovss.n1644 iovss.n1596 9.0005
R7401 iovss.n1644 iovss.n1553 9.0005
R7402 iovss.n1644 iovss.n1598 9.0005
R7403 iovss.n1644 iovss.n1552 9.0005
R7404 iovss.n1644 iovss.n1599 9.0005
R7405 iovss.n1644 iovss.n1551 9.0005
R7406 iovss.n2396 iovss.n1644 9.0005
R7407 iovss.n2394 iovss.n1644 9.0005
R7408 iovss.n1606 iovss.n1569 9.0005
R7409 iovss.n1606 iovss.n1567 9.0005
R7410 iovss.n1606 iovss.n1571 9.0005
R7411 iovss.n1606 iovss.n1566 9.0005
R7412 iovss.n1606 iovss.n1573 9.0005
R7413 iovss.n1606 iovss.n1565 9.0005
R7414 iovss.n1606 iovss.n1575 9.0005
R7415 iovss.n1606 iovss.n1564 9.0005
R7416 iovss.n1606 iovss.n1577 9.0005
R7417 iovss.n1606 iovss.n1563 9.0005
R7418 iovss.n1606 iovss.n1579 9.0005
R7419 iovss.n1606 iovss.n1562 9.0005
R7420 iovss.n1606 iovss.n1581 9.0005
R7421 iovss.n1606 iovss.n1561 9.0005
R7422 iovss.n1606 iovss.n1583 9.0005
R7423 iovss.n1606 iovss.n1560 9.0005
R7424 iovss.n1606 iovss.n1585 9.0005
R7425 iovss.n1606 iovss.n1559 9.0005
R7426 iovss.n1606 iovss.n1587 9.0005
R7427 iovss.n1606 iovss.n1558 9.0005
R7428 iovss.n1606 iovss.n1589 9.0005
R7429 iovss.n1606 iovss.n1557 9.0005
R7430 iovss.n1606 iovss.n1591 9.0005
R7431 iovss.n1606 iovss.n1556 9.0005
R7432 iovss.n1606 iovss.n1593 9.0005
R7433 iovss.n1606 iovss.n1555 9.0005
R7434 iovss.n1606 iovss.n1595 9.0005
R7435 iovss.n1606 iovss.n1554 9.0005
R7436 iovss.n1606 iovss.n1596 9.0005
R7437 iovss.n1606 iovss.n1553 9.0005
R7438 iovss.n1606 iovss.n1598 9.0005
R7439 iovss.n1606 iovss.n1552 9.0005
R7440 iovss.n1606 iovss.n1599 9.0005
R7441 iovss.n1606 iovss.n1551 9.0005
R7442 iovss.n2396 iovss.n1606 9.0005
R7443 iovss.n2394 iovss.n1606 9.0005
R7444 iovss.n1645 iovss.n1569 9.0005
R7445 iovss.n1645 iovss.n1567 9.0005
R7446 iovss.n1645 iovss.n1571 9.0005
R7447 iovss.n1645 iovss.n1566 9.0005
R7448 iovss.n1645 iovss.n1573 9.0005
R7449 iovss.n1645 iovss.n1565 9.0005
R7450 iovss.n1645 iovss.n1575 9.0005
R7451 iovss.n1645 iovss.n1564 9.0005
R7452 iovss.n1645 iovss.n1577 9.0005
R7453 iovss.n1645 iovss.n1563 9.0005
R7454 iovss.n1645 iovss.n1579 9.0005
R7455 iovss.n1645 iovss.n1562 9.0005
R7456 iovss.n1645 iovss.n1581 9.0005
R7457 iovss.n1645 iovss.n1561 9.0005
R7458 iovss.n1645 iovss.n1583 9.0005
R7459 iovss.n1645 iovss.n1560 9.0005
R7460 iovss.n1645 iovss.n1585 9.0005
R7461 iovss.n1645 iovss.n1559 9.0005
R7462 iovss.n1645 iovss.n1587 9.0005
R7463 iovss.n1645 iovss.n1558 9.0005
R7464 iovss.n1645 iovss.n1589 9.0005
R7465 iovss.n1645 iovss.n1557 9.0005
R7466 iovss.n1645 iovss.n1591 9.0005
R7467 iovss.n1645 iovss.n1556 9.0005
R7468 iovss.n1645 iovss.n1593 9.0005
R7469 iovss.n1645 iovss.n1555 9.0005
R7470 iovss.n1645 iovss.n1595 9.0005
R7471 iovss.n1645 iovss.n1554 9.0005
R7472 iovss.n1645 iovss.n1596 9.0005
R7473 iovss.n1645 iovss.n1553 9.0005
R7474 iovss.n1645 iovss.n1598 9.0005
R7475 iovss.n1645 iovss.n1552 9.0005
R7476 iovss.n1645 iovss.n1599 9.0005
R7477 iovss.n1645 iovss.n1551 9.0005
R7478 iovss.n2396 iovss.n1645 9.0005
R7479 iovss.n2394 iovss.n1645 9.0005
R7480 iovss.n1605 iovss.n1569 9.0005
R7481 iovss.n1605 iovss.n1567 9.0005
R7482 iovss.n1605 iovss.n1571 9.0005
R7483 iovss.n1605 iovss.n1566 9.0005
R7484 iovss.n1605 iovss.n1573 9.0005
R7485 iovss.n1605 iovss.n1565 9.0005
R7486 iovss.n1605 iovss.n1575 9.0005
R7487 iovss.n1605 iovss.n1564 9.0005
R7488 iovss.n1605 iovss.n1577 9.0005
R7489 iovss.n1605 iovss.n1563 9.0005
R7490 iovss.n1605 iovss.n1579 9.0005
R7491 iovss.n1605 iovss.n1562 9.0005
R7492 iovss.n1605 iovss.n1581 9.0005
R7493 iovss.n1605 iovss.n1561 9.0005
R7494 iovss.n1605 iovss.n1583 9.0005
R7495 iovss.n1605 iovss.n1560 9.0005
R7496 iovss.n1605 iovss.n1585 9.0005
R7497 iovss.n1605 iovss.n1559 9.0005
R7498 iovss.n1605 iovss.n1587 9.0005
R7499 iovss.n1605 iovss.n1558 9.0005
R7500 iovss.n1605 iovss.n1589 9.0005
R7501 iovss.n1605 iovss.n1557 9.0005
R7502 iovss.n1605 iovss.n1591 9.0005
R7503 iovss.n1605 iovss.n1556 9.0005
R7504 iovss.n1605 iovss.n1593 9.0005
R7505 iovss.n1605 iovss.n1555 9.0005
R7506 iovss.n1605 iovss.n1595 9.0005
R7507 iovss.n1605 iovss.n1554 9.0005
R7508 iovss.n1605 iovss.n1596 9.0005
R7509 iovss.n1605 iovss.n1553 9.0005
R7510 iovss.n1605 iovss.n1598 9.0005
R7511 iovss.n1605 iovss.n1552 9.0005
R7512 iovss.n1605 iovss.n1599 9.0005
R7513 iovss.n1605 iovss.n1551 9.0005
R7514 iovss.n2396 iovss.n1605 9.0005
R7515 iovss.n2394 iovss.n1605 9.0005
R7516 iovss.n1646 iovss.n1569 9.0005
R7517 iovss.n1646 iovss.n1567 9.0005
R7518 iovss.n1646 iovss.n1571 9.0005
R7519 iovss.n1646 iovss.n1566 9.0005
R7520 iovss.n1646 iovss.n1573 9.0005
R7521 iovss.n1646 iovss.n1565 9.0005
R7522 iovss.n1646 iovss.n1575 9.0005
R7523 iovss.n1646 iovss.n1564 9.0005
R7524 iovss.n1646 iovss.n1577 9.0005
R7525 iovss.n1646 iovss.n1563 9.0005
R7526 iovss.n1646 iovss.n1579 9.0005
R7527 iovss.n1646 iovss.n1562 9.0005
R7528 iovss.n1646 iovss.n1581 9.0005
R7529 iovss.n1646 iovss.n1561 9.0005
R7530 iovss.n1646 iovss.n1583 9.0005
R7531 iovss.n1646 iovss.n1560 9.0005
R7532 iovss.n1646 iovss.n1585 9.0005
R7533 iovss.n1646 iovss.n1559 9.0005
R7534 iovss.n1646 iovss.n1587 9.0005
R7535 iovss.n1646 iovss.n1558 9.0005
R7536 iovss.n1646 iovss.n1589 9.0005
R7537 iovss.n1646 iovss.n1557 9.0005
R7538 iovss.n1646 iovss.n1591 9.0005
R7539 iovss.n1646 iovss.n1556 9.0005
R7540 iovss.n1646 iovss.n1593 9.0005
R7541 iovss.n1646 iovss.n1555 9.0005
R7542 iovss.n1646 iovss.n1595 9.0005
R7543 iovss.n1646 iovss.n1554 9.0005
R7544 iovss.n1646 iovss.n1596 9.0005
R7545 iovss.n1646 iovss.n1553 9.0005
R7546 iovss.n1646 iovss.n1598 9.0005
R7547 iovss.n1646 iovss.n1552 9.0005
R7548 iovss.n1646 iovss.n1599 9.0005
R7549 iovss.n1646 iovss.n1551 9.0005
R7550 iovss.n2396 iovss.n1646 9.0005
R7551 iovss.n2394 iovss.n1646 9.0005
R7552 iovss.n1604 iovss.n1569 9.0005
R7553 iovss.n1604 iovss.n1567 9.0005
R7554 iovss.n1604 iovss.n1571 9.0005
R7555 iovss.n1604 iovss.n1566 9.0005
R7556 iovss.n1604 iovss.n1573 9.0005
R7557 iovss.n1604 iovss.n1565 9.0005
R7558 iovss.n1604 iovss.n1575 9.0005
R7559 iovss.n1604 iovss.n1564 9.0005
R7560 iovss.n1604 iovss.n1577 9.0005
R7561 iovss.n1604 iovss.n1563 9.0005
R7562 iovss.n1604 iovss.n1579 9.0005
R7563 iovss.n1604 iovss.n1562 9.0005
R7564 iovss.n1604 iovss.n1581 9.0005
R7565 iovss.n1604 iovss.n1561 9.0005
R7566 iovss.n1604 iovss.n1583 9.0005
R7567 iovss.n1604 iovss.n1560 9.0005
R7568 iovss.n1604 iovss.n1585 9.0005
R7569 iovss.n1604 iovss.n1559 9.0005
R7570 iovss.n1604 iovss.n1587 9.0005
R7571 iovss.n1604 iovss.n1558 9.0005
R7572 iovss.n1604 iovss.n1589 9.0005
R7573 iovss.n1604 iovss.n1557 9.0005
R7574 iovss.n1604 iovss.n1591 9.0005
R7575 iovss.n1604 iovss.n1556 9.0005
R7576 iovss.n1604 iovss.n1593 9.0005
R7577 iovss.n1604 iovss.n1555 9.0005
R7578 iovss.n1604 iovss.n1595 9.0005
R7579 iovss.n1604 iovss.n1554 9.0005
R7580 iovss.n1604 iovss.n1596 9.0005
R7581 iovss.n1604 iovss.n1553 9.0005
R7582 iovss.n1604 iovss.n1598 9.0005
R7583 iovss.n1604 iovss.n1552 9.0005
R7584 iovss.n1604 iovss.n1599 9.0005
R7585 iovss.n1604 iovss.n1551 9.0005
R7586 iovss.n2396 iovss.n1604 9.0005
R7587 iovss.n2394 iovss.n1604 9.0005
R7588 iovss.n1647 iovss.n1569 9.0005
R7589 iovss.n1647 iovss.n1567 9.0005
R7590 iovss.n1647 iovss.n1571 9.0005
R7591 iovss.n1647 iovss.n1566 9.0005
R7592 iovss.n1647 iovss.n1573 9.0005
R7593 iovss.n1647 iovss.n1565 9.0005
R7594 iovss.n1647 iovss.n1575 9.0005
R7595 iovss.n1647 iovss.n1564 9.0005
R7596 iovss.n1647 iovss.n1577 9.0005
R7597 iovss.n1647 iovss.n1563 9.0005
R7598 iovss.n1647 iovss.n1579 9.0005
R7599 iovss.n1647 iovss.n1562 9.0005
R7600 iovss.n1647 iovss.n1581 9.0005
R7601 iovss.n1647 iovss.n1561 9.0005
R7602 iovss.n1647 iovss.n1583 9.0005
R7603 iovss.n1647 iovss.n1560 9.0005
R7604 iovss.n1647 iovss.n1585 9.0005
R7605 iovss.n1647 iovss.n1559 9.0005
R7606 iovss.n1647 iovss.n1587 9.0005
R7607 iovss.n1647 iovss.n1558 9.0005
R7608 iovss.n1647 iovss.n1589 9.0005
R7609 iovss.n1647 iovss.n1557 9.0005
R7610 iovss.n1647 iovss.n1591 9.0005
R7611 iovss.n1647 iovss.n1556 9.0005
R7612 iovss.n1647 iovss.n1593 9.0005
R7613 iovss.n1647 iovss.n1555 9.0005
R7614 iovss.n1647 iovss.n1595 9.0005
R7615 iovss.n1647 iovss.n1554 9.0005
R7616 iovss.n1647 iovss.n1596 9.0005
R7617 iovss.n1647 iovss.n1553 9.0005
R7618 iovss.n1647 iovss.n1598 9.0005
R7619 iovss.n1647 iovss.n1552 9.0005
R7620 iovss.n1647 iovss.n1599 9.0005
R7621 iovss.n1647 iovss.n1551 9.0005
R7622 iovss.n2396 iovss.n1647 9.0005
R7623 iovss.n2394 iovss.n1647 9.0005
R7624 iovss.n1603 iovss.n1569 9.0005
R7625 iovss.n1603 iovss.n1567 9.0005
R7626 iovss.n1603 iovss.n1571 9.0005
R7627 iovss.n1603 iovss.n1566 9.0005
R7628 iovss.n1603 iovss.n1573 9.0005
R7629 iovss.n1603 iovss.n1565 9.0005
R7630 iovss.n1603 iovss.n1575 9.0005
R7631 iovss.n1603 iovss.n1564 9.0005
R7632 iovss.n1603 iovss.n1577 9.0005
R7633 iovss.n1603 iovss.n1563 9.0005
R7634 iovss.n1603 iovss.n1579 9.0005
R7635 iovss.n1603 iovss.n1562 9.0005
R7636 iovss.n1603 iovss.n1581 9.0005
R7637 iovss.n1603 iovss.n1561 9.0005
R7638 iovss.n1603 iovss.n1583 9.0005
R7639 iovss.n1603 iovss.n1560 9.0005
R7640 iovss.n1603 iovss.n1585 9.0005
R7641 iovss.n1603 iovss.n1559 9.0005
R7642 iovss.n1603 iovss.n1587 9.0005
R7643 iovss.n1603 iovss.n1558 9.0005
R7644 iovss.n1603 iovss.n1589 9.0005
R7645 iovss.n1603 iovss.n1557 9.0005
R7646 iovss.n1603 iovss.n1591 9.0005
R7647 iovss.n1603 iovss.n1556 9.0005
R7648 iovss.n1603 iovss.n1593 9.0005
R7649 iovss.n1603 iovss.n1555 9.0005
R7650 iovss.n1603 iovss.n1595 9.0005
R7651 iovss.n1603 iovss.n1554 9.0005
R7652 iovss.n1603 iovss.n1596 9.0005
R7653 iovss.n1603 iovss.n1553 9.0005
R7654 iovss.n1603 iovss.n1598 9.0005
R7655 iovss.n1603 iovss.n1552 9.0005
R7656 iovss.n1603 iovss.n1599 9.0005
R7657 iovss.n1603 iovss.n1551 9.0005
R7658 iovss.n2396 iovss.n1603 9.0005
R7659 iovss.n2394 iovss.n1603 9.0005
R7660 iovss.n1648 iovss.n1569 9.0005
R7661 iovss.n1648 iovss.n1567 9.0005
R7662 iovss.n1648 iovss.n1571 9.0005
R7663 iovss.n1648 iovss.n1566 9.0005
R7664 iovss.n1648 iovss.n1573 9.0005
R7665 iovss.n1648 iovss.n1565 9.0005
R7666 iovss.n1648 iovss.n1575 9.0005
R7667 iovss.n1648 iovss.n1564 9.0005
R7668 iovss.n1648 iovss.n1577 9.0005
R7669 iovss.n1648 iovss.n1563 9.0005
R7670 iovss.n1648 iovss.n1579 9.0005
R7671 iovss.n1648 iovss.n1562 9.0005
R7672 iovss.n1648 iovss.n1581 9.0005
R7673 iovss.n1648 iovss.n1561 9.0005
R7674 iovss.n1648 iovss.n1583 9.0005
R7675 iovss.n1648 iovss.n1560 9.0005
R7676 iovss.n1648 iovss.n1585 9.0005
R7677 iovss.n1648 iovss.n1559 9.0005
R7678 iovss.n1648 iovss.n1587 9.0005
R7679 iovss.n1648 iovss.n1558 9.0005
R7680 iovss.n1648 iovss.n1589 9.0005
R7681 iovss.n1648 iovss.n1557 9.0005
R7682 iovss.n1648 iovss.n1591 9.0005
R7683 iovss.n1648 iovss.n1556 9.0005
R7684 iovss.n1648 iovss.n1593 9.0005
R7685 iovss.n1648 iovss.n1555 9.0005
R7686 iovss.n1648 iovss.n1595 9.0005
R7687 iovss.n1648 iovss.n1554 9.0005
R7688 iovss.n1648 iovss.n1596 9.0005
R7689 iovss.n1648 iovss.n1553 9.0005
R7690 iovss.n1648 iovss.n1598 9.0005
R7691 iovss.n1648 iovss.n1552 9.0005
R7692 iovss.n1648 iovss.n1599 9.0005
R7693 iovss.n1648 iovss.n1551 9.0005
R7694 iovss.n2396 iovss.n1648 9.0005
R7695 iovss.n2394 iovss.n1648 9.0005
R7696 iovss.n1602 iovss.n1569 9.0005
R7697 iovss.n1602 iovss.n1567 9.0005
R7698 iovss.n1602 iovss.n1571 9.0005
R7699 iovss.n1602 iovss.n1566 9.0005
R7700 iovss.n1602 iovss.n1573 9.0005
R7701 iovss.n1602 iovss.n1565 9.0005
R7702 iovss.n1602 iovss.n1575 9.0005
R7703 iovss.n1602 iovss.n1564 9.0005
R7704 iovss.n1602 iovss.n1577 9.0005
R7705 iovss.n1602 iovss.n1563 9.0005
R7706 iovss.n1602 iovss.n1579 9.0005
R7707 iovss.n1602 iovss.n1562 9.0005
R7708 iovss.n1602 iovss.n1581 9.0005
R7709 iovss.n1602 iovss.n1561 9.0005
R7710 iovss.n1602 iovss.n1583 9.0005
R7711 iovss.n1602 iovss.n1560 9.0005
R7712 iovss.n1602 iovss.n1585 9.0005
R7713 iovss.n1602 iovss.n1559 9.0005
R7714 iovss.n1602 iovss.n1587 9.0005
R7715 iovss.n1602 iovss.n1558 9.0005
R7716 iovss.n1602 iovss.n1589 9.0005
R7717 iovss.n1602 iovss.n1557 9.0005
R7718 iovss.n1602 iovss.n1591 9.0005
R7719 iovss.n1602 iovss.n1556 9.0005
R7720 iovss.n1602 iovss.n1593 9.0005
R7721 iovss.n1602 iovss.n1555 9.0005
R7722 iovss.n1602 iovss.n1595 9.0005
R7723 iovss.n1602 iovss.n1554 9.0005
R7724 iovss.n1602 iovss.n1596 9.0005
R7725 iovss.n1602 iovss.n1553 9.0005
R7726 iovss.n1602 iovss.n1598 9.0005
R7727 iovss.n1602 iovss.n1552 9.0005
R7728 iovss.n1602 iovss.n1599 9.0005
R7729 iovss.n1602 iovss.n1551 9.0005
R7730 iovss.n2396 iovss.n1602 9.0005
R7731 iovss.n2394 iovss.n1602 9.0005
R7732 iovss.n1649 iovss.n1569 9.0005
R7733 iovss.n1649 iovss.n1567 9.0005
R7734 iovss.n1649 iovss.n1571 9.0005
R7735 iovss.n1649 iovss.n1566 9.0005
R7736 iovss.n1649 iovss.n1573 9.0005
R7737 iovss.n1649 iovss.n1565 9.0005
R7738 iovss.n1649 iovss.n1575 9.0005
R7739 iovss.n1649 iovss.n1564 9.0005
R7740 iovss.n1649 iovss.n1577 9.0005
R7741 iovss.n1649 iovss.n1563 9.0005
R7742 iovss.n1649 iovss.n1579 9.0005
R7743 iovss.n1649 iovss.n1562 9.0005
R7744 iovss.n1649 iovss.n1581 9.0005
R7745 iovss.n1649 iovss.n1561 9.0005
R7746 iovss.n1649 iovss.n1583 9.0005
R7747 iovss.n1649 iovss.n1560 9.0005
R7748 iovss.n1649 iovss.n1585 9.0005
R7749 iovss.n1649 iovss.n1559 9.0005
R7750 iovss.n1649 iovss.n1587 9.0005
R7751 iovss.n1649 iovss.n1558 9.0005
R7752 iovss.n1649 iovss.n1589 9.0005
R7753 iovss.n1649 iovss.n1557 9.0005
R7754 iovss.n1649 iovss.n1591 9.0005
R7755 iovss.n1649 iovss.n1556 9.0005
R7756 iovss.n1649 iovss.n1593 9.0005
R7757 iovss.n1649 iovss.n1555 9.0005
R7758 iovss.n1649 iovss.n1595 9.0005
R7759 iovss.n1649 iovss.n1554 9.0005
R7760 iovss.n1649 iovss.n1596 9.0005
R7761 iovss.n1649 iovss.n1553 9.0005
R7762 iovss.n1649 iovss.n1598 9.0005
R7763 iovss.n1649 iovss.n1552 9.0005
R7764 iovss.n1649 iovss.n1599 9.0005
R7765 iovss.n1649 iovss.n1551 9.0005
R7766 iovss.n2396 iovss.n1649 9.0005
R7767 iovss.n2394 iovss.n1649 9.0005
R7768 iovss.n1601 iovss.n1569 9.0005
R7769 iovss.n1601 iovss.n1567 9.0005
R7770 iovss.n1601 iovss.n1571 9.0005
R7771 iovss.n1601 iovss.n1566 9.0005
R7772 iovss.n1601 iovss.n1573 9.0005
R7773 iovss.n1601 iovss.n1565 9.0005
R7774 iovss.n1601 iovss.n1575 9.0005
R7775 iovss.n1601 iovss.n1564 9.0005
R7776 iovss.n1601 iovss.n1577 9.0005
R7777 iovss.n1601 iovss.n1563 9.0005
R7778 iovss.n1601 iovss.n1579 9.0005
R7779 iovss.n1601 iovss.n1562 9.0005
R7780 iovss.n1601 iovss.n1581 9.0005
R7781 iovss.n1601 iovss.n1561 9.0005
R7782 iovss.n1601 iovss.n1583 9.0005
R7783 iovss.n1601 iovss.n1560 9.0005
R7784 iovss.n1601 iovss.n1585 9.0005
R7785 iovss.n1601 iovss.n1559 9.0005
R7786 iovss.n1601 iovss.n1587 9.0005
R7787 iovss.n1601 iovss.n1558 9.0005
R7788 iovss.n1601 iovss.n1589 9.0005
R7789 iovss.n1601 iovss.n1557 9.0005
R7790 iovss.n1601 iovss.n1591 9.0005
R7791 iovss.n1601 iovss.n1556 9.0005
R7792 iovss.n1601 iovss.n1593 9.0005
R7793 iovss.n1601 iovss.n1555 9.0005
R7794 iovss.n1601 iovss.n1595 9.0005
R7795 iovss.n1601 iovss.n1554 9.0005
R7796 iovss.n1601 iovss.n1596 9.0005
R7797 iovss.n1601 iovss.n1553 9.0005
R7798 iovss.n1601 iovss.n1598 9.0005
R7799 iovss.n1601 iovss.n1552 9.0005
R7800 iovss.n1601 iovss.n1599 9.0005
R7801 iovss.n1601 iovss.n1551 9.0005
R7802 iovss.n2396 iovss.n1601 9.0005
R7803 iovss.n2394 iovss.n1601 9.0005
R7804 iovss.n2395 iovss.n1569 9.0005
R7805 iovss.n2395 iovss.n1567 9.0005
R7806 iovss.n2395 iovss.n1571 9.0005
R7807 iovss.n2395 iovss.n1566 9.0005
R7808 iovss.n2395 iovss.n1573 9.0005
R7809 iovss.n2395 iovss.n1565 9.0005
R7810 iovss.n2395 iovss.n1575 9.0005
R7811 iovss.n2395 iovss.n1564 9.0005
R7812 iovss.n2395 iovss.n1577 9.0005
R7813 iovss.n2395 iovss.n1563 9.0005
R7814 iovss.n2395 iovss.n1579 9.0005
R7815 iovss.n2395 iovss.n1562 9.0005
R7816 iovss.n2395 iovss.n1581 9.0005
R7817 iovss.n2395 iovss.n1561 9.0005
R7818 iovss.n2395 iovss.n1583 9.0005
R7819 iovss.n2395 iovss.n1560 9.0005
R7820 iovss.n2395 iovss.n1585 9.0005
R7821 iovss.n2395 iovss.n1559 9.0005
R7822 iovss.n2395 iovss.n1587 9.0005
R7823 iovss.n2395 iovss.n1558 9.0005
R7824 iovss.n2395 iovss.n1589 9.0005
R7825 iovss.n2395 iovss.n1557 9.0005
R7826 iovss.n2395 iovss.n1591 9.0005
R7827 iovss.n2395 iovss.n1556 9.0005
R7828 iovss.n2395 iovss.n1593 9.0005
R7829 iovss.n2395 iovss.n1555 9.0005
R7830 iovss.n2395 iovss.n1595 9.0005
R7831 iovss.n2395 iovss.n1554 9.0005
R7832 iovss.n2395 iovss.n1596 9.0005
R7833 iovss.n2395 iovss.n1553 9.0005
R7834 iovss.n2395 iovss.n1598 9.0005
R7835 iovss.n2395 iovss.n1552 9.0005
R7836 iovss.n2395 iovss.n1599 9.0005
R7837 iovss.n2395 iovss.n1551 9.0005
R7838 iovss.n2396 iovss.n2395 9.0005
R7839 iovss.n2395 iovss.n2394 9.0005
R7840 iovss.n1600 iovss.n1569 9.0005
R7841 iovss.n1600 iovss.n1567 9.0005
R7842 iovss.n1600 iovss.n1571 9.0005
R7843 iovss.n1600 iovss.n1566 9.0005
R7844 iovss.n1600 iovss.n1573 9.0005
R7845 iovss.n1600 iovss.n1565 9.0005
R7846 iovss.n1600 iovss.n1575 9.0005
R7847 iovss.n1600 iovss.n1564 9.0005
R7848 iovss.n1600 iovss.n1577 9.0005
R7849 iovss.n1600 iovss.n1563 9.0005
R7850 iovss.n1600 iovss.n1579 9.0005
R7851 iovss.n1600 iovss.n1562 9.0005
R7852 iovss.n1600 iovss.n1581 9.0005
R7853 iovss.n1600 iovss.n1561 9.0005
R7854 iovss.n1600 iovss.n1583 9.0005
R7855 iovss.n1600 iovss.n1560 9.0005
R7856 iovss.n1600 iovss.n1585 9.0005
R7857 iovss.n1600 iovss.n1559 9.0005
R7858 iovss.n1600 iovss.n1587 9.0005
R7859 iovss.n1600 iovss.n1558 9.0005
R7860 iovss.n1600 iovss.n1589 9.0005
R7861 iovss.n1600 iovss.n1557 9.0005
R7862 iovss.n1600 iovss.n1591 9.0005
R7863 iovss.n1600 iovss.n1556 9.0005
R7864 iovss.n1600 iovss.n1593 9.0005
R7865 iovss.n1600 iovss.n1555 9.0005
R7866 iovss.n1600 iovss.n1595 9.0005
R7867 iovss.n1600 iovss.n1554 9.0005
R7868 iovss.n1600 iovss.n1596 9.0005
R7869 iovss.n1600 iovss.n1553 9.0005
R7870 iovss.n1600 iovss.n1598 9.0005
R7871 iovss.n1600 iovss.n1552 9.0005
R7872 iovss.n1600 iovss.n1599 9.0005
R7873 iovss.n1600 iovss.n1551 9.0005
R7874 iovss.n2396 iovss.n1600 9.0005
R7875 iovss.n2394 iovss.n1600 9.0005
R7876 iovss.n2397 iovss.n1569 9.0005
R7877 iovss.n2397 iovss.n1567 9.0005
R7878 iovss.n2397 iovss.n1571 9.0005
R7879 iovss.n2397 iovss.n1566 9.0005
R7880 iovss.n2397 iovss.n1573 9.0005
R7881 iovss.n2397 iovss.n1565 9.0005
R7882 iovss.n2397 iovss.n1575 9.0005
R7883 iovss.n2397 iovss.n1564 9.0005
R7884 iovss.n2397 iovss.n1577 9.0005
R7885 iovss.n2397 iovss.n1563 9.0005
R7886 iovss.n2397 iovss.n1579 9.0005
R7887 iovss.n2397 iovss.n1562 9.0005
R7888 iovss.n2397 iovss.n1581 9.0005
R7889 iovss.n2397 iovss.n1561 9.0005
R7890 iovss.n2397 iovss.n1583 9.0005
R7891 iovss.n2397 iovss.n1560 9.0005
R7892 iovss.n2397 iovss.n1585 9.0005
R7893 iovss.n2397 iovss.n1559 9.0005
R7894 iovss.n2397 iovss.n1587 9.0005
R7895 iovss.n2397 iovss.n1558 9.0005
R7896 iovss.n2397 iovss.n1589 9.0005
R7897 iovss.n2397 iovss.n1557 9.0005
R7898 iovss.n2397 iovss.n1591 9.0005
R7899 iovss.n2397 iovss.n1556 9.0005
R7900 iovss.n2397 iovss.n1593 9.0005
R7901 iovss.n2397 iovss.n1555 9.0005
R7902 iovss.n2397 iovss.n1595 9.0005
R7903 iovss.n2397 iovss.n1554 9.0005
R7904 iovss.n2397 iovss.n1596 9.0005
R7905 iovss.n2397 iovss.n1553 9.0005
R7906 iovss.n2397 iovss.n1598 9.0005
R7907 iovss.n2397 iovss.n1552 9.0005
R7908 iovss.n2397 iovss.n1599 9.0005
R7909 iovss.n2397 iovss.n1551 9.0005
R7910 iovss.n2397 iovss.n2396 9.0005
R7911 iovss.n2452 iovss.n2398 9.0005
R7912 iovss.n2454 iovss.n2398 9.0005
R7913 iovss.n2460 iovss.n2398 9.0005
R7914 iovss.n2451 iovss.n2398 9.0005
R7915 iovss.n2445 iovss.n2398 9.0005
R7916 iovss.n2443 iovss.n2398 9.0005
R7917 iovss.n2427 iovss.n2398 9.0005
R7918 iovss.n2470 iovss.n2398 9.0005
R7919 iovss.n2476 iovss.n2398 9.0005
R7920 iovss.n2478 iovss.n2398 9.0005
R7921 iovss.n2484 iovss.n2398 9.0005
R7922 iovss.n2426 iovss.n2398 9.0005
R7923 iovss.n2420 iovss.n2398 9.0005
R7924 iovss.n2418 iovss.n2398 9.0005
R7925 iovss.n2403 iovss.n2398 9.0005
R7926 iovss.n2494 iovss.n2398 9.0005
R7927 iovss.n2500 iovss.n2398 9.0005
R7928 iovss.n2510 iovss.n2398 9.0005
R7929 iovss.n2452 iovss.n2399 9.0005
R7930 iovss.n2505 iovss.n2399 9.0005
R7931 iovss.n2510 iovss.n2399 9.0005
R7932 iovss.n2452 iovss.n1444 9.0005
R7933 iovss.n2454 iovss.n1444 9.0005
R7934 iovss.n2456 iovss.n1444 9.0005
R7935 iovss.n2458 iovss.n1444 9.0005
R7936 iovss.n2460 iovss.n1444 9.0005
R7937 iovss.n2451 iovss.n1444 9.0005
R7938 iovss.n2449 iovss.n1444 9.0005
R7939 iovss.n2447 iovss.n1444 9.0005
R7940 iovss.n2445 iovss.n1444 9.0005
R7941 iovss.n2443 iovss.n1444 9.0005
R7942 iovss.n2441 iovss.n1444 9.0005
R7943 iovss.n2439 iovss.n1444 9.0005
R7944 iovss.n2427 iovss.n1444 9.0005
R7945 iovss.n2470 iovss.n1444 9.0005
R7946 iovss.n2472 iovss.n1444 9.0005
R7947 iovss.n2474 iovss.n1444 9.0005
R7948 iovss.n2476 iovss.n1444 9.0005
R7949 iovss.n2478 iovss.n1444 9.0005
R7950 iovss.n2480 iovss.n1444 9.0005
R7951 iovss.n2482 iovss.n1444 9.0005
R7952 iovss.n2484 iovss.n1444 9.0005
R7953 iovss.n2426 iovss.n1444 9.0005
R7954 iovss.n2424 iovss.n1444 9.0005
R7955 iovss.n2422 iovss.n1444 9.0005
R7956 iovss.n2420 iovss.n1444 9.0005
R7957 iovss.n2418 iovss.n1444 9.0005
R7958 iovss.n2416 iovss.n1444 9.0005
R7959 iovss.n2414 iovss.n1444 9.0005
R7960 iovss.n2403 iovss.n1444 9.0005
R7961 iovss.n2494 iovss.n1444 9.0005
R7962 iovss.n2496 iovss.n1444 9.0005
R7963 iovss.n2498 iovss.n1444 9.0005
R7964 iovss.n2500 iovss.n1444 9.0005
R7965 iovss.n2510 iovss.n1444 9.0005
R7966 iovss.n2452 iovss.n1443 9.0005
R7967 iovss.n2454 iovss.n1443 9.0005
R7968 iovss.n2456 iovss.n1443 9.0005
R7969 iovss.n2458 iovss.n1443 9.0005
R7970 iovss.n2460 iovss.n1443 9.0005
R7971 iovss.n2451 iovss.n1443 9.0005
R7972 iovss.n2449 iovss.n1443 9.0005
R7973 iovss.n2447 iovss.n1443 9.0005
R7974 iovss.n2445 iovss.n1443 9.0005
R7975 iovss.n2443 iovss.n1443 9.0005
R7976 iovss.n2441 iovss.n1443 9.0005
R7977 iovss.n2439 iovss.n1443 9.0005
R7978 iovss.n2427 iovss.n1443 9.0005
R7979 iovss.n2470 iovss.n1443 9.0005
R7980 iovss.n2472 iovss.n1443 9.0005
R7981 iovss.n2474 iovss.n1443 9.0005
R7982 iovss.n2476 iovss.n1443 9.0005
R7983 iovss.n2478 iovss.n1443 9.0005
R7984 iovss.n2480 iovss.n1443 9.0005
R7985 iovss.n2482 iovss.n1443 9.0005
R7986 iovss.n2484 iovss.n1443 9.0005
R7987 iovss.n2426 iovss.n1443 9.0005
R7988 iovss.n2424 iovss.n1443 9.0005
R7989 iovss.n2422 iovss.n1443 9.0005
R7990 iovss.n2420 iovss.n1443 9.0005
R7991 iovss.n2418 iovss.n1443 9.0005
R7992 iovss.n2416 iovss.n1443 9.0005
R7993 iovss.n2414 iovss.n1443 9.0005
R7994 iovss.n2403 iovss.n1443 9.0005
R7995 iovss.n2494 iovss.n1443 9.0005
R7996 iovss.n2496 iovss.n1443 9.0005
R7997 iovss.n2498 iovss.n1443 9.0005
R7998 iovss.n2500 iovss.n1443 9.0005
R7999 iovss.n2503 iovss.n1443 9.0005
R8000 iovss.n2505 iovss.n1443 9.0005
R8001 iovss.n2510 iovss.n1443 9.0005
R8002 iovss.n2452 iovss.n1548 9.0005
R8003 iovss.n2454 iovss.n1548 9.0005
R8004 iovss.n2456 iovss.n1548 9.0005
R8005 iovss.n2458 iovss.n1548 9.0005
R8006 iovss.n2460 iovss.n1548 9.0005
R8007 iovss.n2451 iovss.n1548 9.0005
R8008 iovss.n2449 iovss.n1548 9.0005
R8009 iovss.n2447 iovss.n1548 9.0005
R8010 iovss.n2445 iovss.n1548 9.0005
R8011 iovss.n2443 iovss.n1548 9.0005
R8012 iovss.n2441 iovss.n1548 9.0005
R8013 iovss.n2439 iovss.n1548 9.0005
R8014 iovss.n2427 iovss.n1548 9.0005
R8015 iovss.n2470 iovss.n1548 9.0005
R8016 iovss.n2472 iovss.n1548 9.0005
R8017 iovss.n2474 iovss.n1548 9.0005
R8018 iovss.n2476 iovss.n1548 9.0005
R8019 iovss.n2478 iovss.n1548 9.0005
R8020 iovss.n2480 iovss.n1548 9.0005
R8021 iovss.n2482 iovss.n1548 9.0005
R8022 iovss.n2484 iovss.n1548 9.0005
R8023 iovss.n2426 iovss.n1548 9.0005
R8024 iovss.n2424 iovss.n1548 9.0005
R8025 iovss.n2422 iovss.n1548 9.0005
R8026 iovss.n2420 iovss.n1548 9.0005
R8027 iovss.n2418 iovss.n1548 9.0005
R8028 iovss.n2416 iovss.n1548 9.0005
R8029 iovss.n2414 iovss.n1548 9.0005
R8030 iovss.n2403 iovss.n1548 9.0005
R8031 iovss.n2494 iovss.n1548 9.0005
R8032 iovss.n2496 iovss.n1548 9.0005
R8033 iovss.n2498 iovss.n1548 9.0005
R8034 iovss.n2500 iovss.n1548 9.0005
R8035 iovss.n2505 iovss.n1548 9.0005
R8036 iovss.n2510 iovss.n1548 9.0005
R8037 iovss.n2452 iovss.n2400 9.0005
R8038 iovss.n2454 iovss.n2400 9.0005
R8039 iovss.n2456 iovss.n2400 9.0005
R8040 iovss.n2458 iovss.n2400 9.0005
R8041 iovss.n2460 iovss.n2400 9.0005
R8042 iovss.n2451 iovss.n2400 9.0005
R8043 iovss.n2449 iovss.n2400 9.0005
R8044 iovss.n2447 iovss.n2400 9.0005
R8045 iovss.n2445 iovss.n2400 9.0005
R8046 iovss.n2443 iovss.n2400 9.0005
R8047 iovss.n2441 iovss.n2400 9.0005
R8048 iovss.n2439 iovss.n2400 9.0005
R8049 iovss.n2427 iovss.n2400 9.0005
R8050 iovss.n2470 iovss.n2400 9.0005
R8051 iovss.n2472 iovss.n2400 9.0005
R8052 iovss.n2474 iovss.n2400 9.0005
R8053 iovss.n2476 iovss.n2400 9.0005
R8054 iovss.n2478 iovss.n2400 9.0005
R8055 iovss.n2480 iovss.n2400 9.0005
R8056 iovss.n2482 iovss.n2400 9.0005
R8057 iovss.n2484 iovss.n2400 9.0005
R8058 iovss.n2426 iovss.n2400 9.0005
R8059 iovss.n2424 iovss.n2400 9.0005
R8060 iovss.n2422 iovss.n2400 9.0005
R8061 iovss.n2420 iovss.n2400 9.0005
R8062 iovss.n2418 iovss.n2400 9.0005
R8063 iovss.n2416 iovss.n2400 9.0005
R8064 iovss.n2414 iovss.n2400 9.0005
R8065 iovss.n2403 iovss.n2400 9.0005
R8066 iovss.n2494 iovss.n2400 9.0005
R8067 iovss.n2496 iovss.n2400 9.0005
R8068 iovss.n2498 iovss.n2400 9.0005
R8069 iovss.n2500 iovss.n2400 9.0005
R8070 iovss.n2505 iovss.n2400 9.0005
R8071 iovss.n2900 iovss.n1225 9.0005
R8072 iovss.n1225 iovss.n1219 9.0005
R8073 iovss.n2789 iovss.n1219 9.0005
R8074 iovss.n2794 iovss.n1219 9.0005
R8075 iovss.n2792 iovss.n1219 9.0005
R8076 iovss.n2799 iovss.n1219 9.0005
R8077 iovss.n2797 iovss.n1219 9.0005
R8078 iovss.n2804 iovss.n1219 9.0005
R8079 iovss.n2802 iovss.n1219 9.0005
R8080 iovss.n2809 iovss.n1219 9.0005
R8081 iovss.n2807 iovss.n1219 9.0005
R8082 iovss.n2814 iovss.n1219 9.0005
R8083 iovss.n2812 iovss.n1219 9.0005
R8084 iovss.n2819 iovss.n1219 9.0005
R8085 iovss.n2817 iovss.n1219 9.0005
R8086 iovss.n2824 iovss.n1219 9.0005
R8087 iovss.n2822 iovss.n1219 9.0005
R8088 iovss.n2829 iovss.n1219 9.0005
R8089 iovss.n2827 iovss.n1219 9.0005
R8090 iovss.n2834 iovss.n1219 9.0005
R8091 iovss.n2832 iovss.n1219 9.0005
R8092 iovss.n2839 iovss.n1219 9.0005
R8093 iovss.n2837 iovss.n1219 9.0005
R8094 iovss.n2844 iovss.n1219 9.0005
R8095 iovss.n2842 iovss.n1219 9.0005
R8096 iovss.n2849 iovss.n1219 9.0005
R8097 iovss.n2847 iovss.n1219 9.0005
R8098 iovss.n2854 iovss.n1219 9.0005
R8099 iovss.n2852 iovss.n1219 9.0005
R8100 iovss.n2859 iovss.n1219 9.0005
R8101 iovss.n2857 iovss.n1219 9.0005
R8102 iovss.n2864 iovss.n1219 9.0005
R8103 iovss.n2862 iovss.n1219 9.0005
R8104 iovss.n2869 iovss.n1219 9.0005
R8105 iovss.n2867 iovss.n1219 9.0005
R8106 iovss.n2874 iovss.n1219 9.0005
R8107 iovss.n2872 iovss.n1219 9.0005
R8108 iovss.n2879 iovss.n1219 9.0005
R8109 iovss.n2877 iovss.n1219 9.0005
R8110 iovss.n2884 iovss.n1219 9.0005
R8111 iovss.n2882 iovss.n1219 9.0005
R8112 iovss.n2887 iovss.n1219 9.0005
R8113 iovss.n2889 iovss.n1219 9.0005
R8114 iovss.n2892 iovss.n1219 9.0005
R8115 iovss.n2900 iovss.n2899 9.0005
R8116 iovss.n2754 iovss.n2602 9.0005
R8117 iovss.n2754 iovss.n2753 9.0005
R8118 iovss.n2753 iovss.n2645 9.0005
R8119 iovss.n2753 iovss.n2648 9.0005
R8120 iovss.n2753 iovss.n2644 9.0005
R8121 iovss.n2753 iovss.n2651 9.0005
R8122 iovss.n2753 iovss.n2642 9.0005
R8123 iovss.n2753 iovss.n2654 9.0005
R8124 iovss.n2753 iovss.n2640 9.0005
R8125 iovss.n2753 iovss.n2657 9.0005
R8126 iovss.n2753 iovss.n2638 9.0005
R8127 iovss.n2753 iovss.n2660 9.0005
R8128 iovss.n2753 iovss.n2636 9.0005
R8129 iovss.n2753 iovss.n2663 9.0005
R8130 iovss.n2753 iovss.n2634 9.0005
R8131 iovss.n2753 iovss.n2666 9.0005
R8132 iovss.n2753 iovss.n2632 9.0005
R8133 iovss.n2753 iovss.n2669 9.0005
R8134 iovss.n2753 iovss.n2630 9.0005
R8135 iovss.n2753 iovss.n2672 9.0005
R8136 iovss.n2753 iovss.n2628 9.0005
R8137 iovss.n2753 iovss.n2675 9.0005
R8138 iovss.n2753 iovss.n2626 9.0005
R8139 iovss.n2753 iovss.n2678 9.0005
R8140 iovss.n2753 iovss.n2624 9.0005
R8141 iovss.n2753 iovss.n2681 9.0005
R8142 iovss.n2753 iovss.n2622 9.0005
R8143 iovss.n2753 iovss.n2684 9.0005
R8144 iovss.n2753 iovss.n2620 9.0005
R8145 iovss.n2753 iovss.n2687 9.0005
R8146 iovss.n2753 iovss.n2618 9.0005
R8147 iovss.n2753 iovss.n2690 9.0005
R8148 iovss.n2753 iovss.n2616 9.0005
R8149 iovss.n2753 iovss.n2693 9.0005
R8150 iovss.n2753 iovss.n2614 9.0005
R8151 iovss.n2753 iovss.n2696 9.0005
R8152 iovss.n2753 iovss.n2612 9.0005
R8153 iovss.n2753 iovss.n2699 9.0005
R8154 iovss.n2753 iovss.n2610 9.0005
R8155 iovss.n2753 iovss.n2702 9.0005
R8156 iovss.n2753 iovss.n2608 9.0005
R8157 iovss.n2753 iovss.n2705 9.0005
R8158 iovss.n2753 iovss.n2606 9.0005
R8159 iovss.n2753 iovss.n2708 9.0005
R8160 iovss.n2753 iovss.n2604 9.0005
R8161 iovss.n1381 iovss.n1340 9.0005
R8162 iovss.n2760 iovss.n1346 9.0005
R8163 iovss.n2760 iovss.n1343 9.0005
R8164 iovss.n2760 iovss.n2759 9.0005
R8165 iovss.n2760 iovss.n1342 9.0005
R8166 iovss.n2761 iovss.n1340 9.0005
R8167 iovss.n2761 iovss.n2760 9.0005
R8168 iovss.n2765 iovss.n1312 9.0005
R8169 iovss.n2773 iovss.n2765 9.0005
R8170 iovss.n2773 iovss.n1318 9.0005
R8171 iovss.n2773 iovss.n2769 9.0005
R8172 iovss.n2773 iovss.n1316 9.0005
R8173 iovss.n2773 iovss.n2772 9.0005
R8174 iovss.n2774 iovss.n2773 9.0005
R8175 iovss.n219 iovss.n172 9.0005
R8176 iovss.n248 iovss.n172 9.0005
R8177 iovss.n205 iovss.n172 9.0005
R8178 iovss.n251 iovss.n172 9.0005
R8179 iovss.n3427 iovss.n172 9.0005
R8180 iovss.n3426 iovss.n219 9.0005
R8181 iovss.n3426 iovss.n222 9.0005
R8182 iovss.n3426 iovss.n217 9.0005
R8183 iovss.n3426 iovss.n226 9.0005
R8184 iovss.n3426 iovss.n215 9.0005
R8185 iovss.n3426 iovss.n230 9.0005
R8186 iovss.n3426 iovss.n213 9.0005
R8187 iovss.n3426 iovss.n234 9.0005
R8188 iovss.n3426 iovss.n211 9.0005
R8189 iovss.n3426 iovss.n237 9.0005
R8190 iovss.n3426 iovss.n210 9.0005
R8191 iovss.n3426 iovss.n241 9.0005
R8192 iovss.n3426 iovss.n253 9.0005
R8193 iovss.n3427 iovss.n3426 9.0005
R8194 iovss.n219 iovss.n184 9.0005
R8195 iovss.n222 iovss.n184 9.0005
R8196 iovss.n218 iovss.n184 9.0005
R8197 iovss.n224 iovss.n184 9.0005
R8198 iovss.n217 iovss.n184 9.0005
R8199 iovss.n226 iovss.n184 9.0005
R8200 iovss.n216 iovss.n184 9.0005
R8201 iovss.n228 iovss.n184 9.0005
R8202 iovss.n215 iovss.n184 9.0005
R8203 iovss.n230 iovss.n184 9.0005
R8204 iovss.n214 iovss.n184 9.0005
R8205 iovss.n232 iovss.n184 9.0005
R8206 iovss.n213 iovss.n184 9.0005
R8207 iovss.n234 iovss.n184 9.0005
R8208 iovss.n212 iovss.n184 9.0005
R8209 iovss.n236 iovss.n184 9.0005
R8210 iovss.n211 iovss.n184 9.0005
R8211 iovss.n237 iovss.n184 9.0005
R8212 iovss.n3429 iovss.n184 9.0005
R8213 iovss.n239 iovss.n184 9.0005
R8214 iovss.n210 iovss.n184 9.0005
R8215 iovss.n241 iovss.n184 9.0005
R8216 iovss.n209 iovss.n184 9.0005
R8217 iovss.n243 iovss.n184 9.0005
R8218 iovss.n208 iovss.n184 9.0005
R8219 iovss.n245 iovss.n184 9.0005
R8220 iovss.n207 iovss.n184 9.0005
R8221 iovss.n247 iovss.n184 9.0005
R8222 iovss.n206 iovss.n184 9.0005
R8223 iovss.n248 iovss.n184 9.0005
R8224 iovss.n205 iovss.n184 9.0005
R8225 iovss.n250 iovss.n184 9.0005
R8226 iovss.n204 iovss.n184 9.0005
R8227 iovss.n251 iovss.n184 9.0005
R8228 iovss.n253 iovss.n184 9.0005
R8229 iovss.n3427 iovss.n184 9.0005
R8230 iovss.n219 iovss.n186 9.0005
R8231 iovss.n222 iovss.n186 9.0005
R8232 iovss.n218 iovss.n186 9.0005
R8233 iovss.n224 iovss.n186 9.0005
R8234 iovss.n217 iovss.n186 9.0005
R8235 iovss.n226 iovss.n186 9.0005
R8236 iovss.n216 iovss.n186 9.0005
R8237 iovss.n228 iovss.n186 9.0005
R8238 iovss.n215 iovss.n186 9.0005
R8239 iovss.n230 iovss.n186 9.0005
R8240 iovss.n214 iovss.n186 9.0005
R8241 iovss.n232 iovss.n186 9.0005
R8242 iovss.n213 iovss.n186 9.0005
R8243 iovss.n234 iovss.n186 9.0005
R8244 iovss.n212 iovss.n186 9.0005
R8245 iovss.n236 iovss.n186 9.0005
R8246 iovss.n211 iovss.n186 9.0005
R8247 iovss.n237 iovss.n186 9.0005
R8248 iovss.n3429 iovss.n186 9.0005
R8249 iovss.n239 iovss.n186 9.0005
R8250 iovss.n210 iovss.n186 9.0005
R8251 iovss.n241 iovss.n186 9.0005
R8252 iovss.n209 iovss.n186 9.0005
R8253 iovss.n243 iovss.n186 9.0005
R8254 iovss.n208 iovss.n186 9.0005
R8255 iovss.n245 iovss.n186 9.0005
R8256 iovss.n207 iovss.n186 9.0005
R8257 iovss.n247 iovss.n186 9.0005
R8258 iovss.n206 iovss.n186 9.0005
R8259 iovss.n248 iovss.n186 9.0005
R8260 iovss.n205 iovss.n186 9.0005
R8261 iovss.n250 iovss.n186 9.0005
R8262 iovss.n204 iovss.n186 9.0005
R8263 iovss.n251 iovss.n186 9.0005
R8264 iovss.n253 iovss.n186 9.0005
R8265 iovss.n3427 iovss.n186 9.0005
R8266 iovss.n219 iovss.n183 9.0005
R8267 iovss.n222 iovss.n183 9.0005
R8268 iovss.n218 iovss.n183 9.0005
R8269 iovss.n224 iovss.n183 9.0005
R8270 iovss.n217 iovss.n183 9.0005
R8271 iovss.n226 iovss.n183 9.0005
R8272 iovss.n216 iovss.n183 9.0005
R8273 iovss.n228 iovss.n183 9.0005
R8274 iovss.n215 iovss.n183 9.0005
R8275 iovss.n230 iovss.n183 9.0005
R8276 iovss.n214 iovss.n183 9.0005
R8277 iovss.n232 iovss.n183 9.0005
R8278 iovss.n213 iovss.n183 9.0005
R8279 iovss.n234 iovss.n183 9.0005
R8280 iovss.n212 iovss.n183 9.0005
R8281 iovss.n236 iovss.n183 9.0005
R8282 iovss.n211 iovss.n183 9.0005
R8283 iovss.n237 iovss.n183 9.0005
R8284 iovss.n3429 iovss.n183 9.0005
R8285 iovss.n239 iovss.n183 9.0005
R8286 iovss.n210 iovss.n183 9.0005
R8287 iovss.n241 iovss.n183 9.0005
R8288 iovss.n209 iovss.n183 9.0005
R8289 iovss.n243 iovss.n183 9.0005
R8290 iovss.n208 iovss.n183 9.0005
R8291 iovss.n245 iovss.n183 9.0005
R8292 iovss.n207 iovss.n183 9.0005
R8293 iovss.n247 iovss.n183 9.0005
R8294 iovss.n206 iovss.n183 9.0005
R8295 iovss.n248 iovss.n183 9.0005
R8296 iovss.n205 iovss.n183 9.0005
R8297 iovss.n250 iovss.n183 9.0005
R8298 iovss.n204 iovss.n183 9.0005
R8299 iovss.n251 iovss.n183 9.0005
R8300 iovss.n253 iovss.n183 9.0005
R8301 iovss.n3427 iovss.n183 9.0005
R8302 iovss.n219 iovss.n187 9.0005
R8303 iovss.n222 iovss.n187 9.0005
R8304 iovss.n218 iovss.n187 9.0005
R8305 iovss.n224 iovss.n187 9.0005
R8306 iovss.n217 iovss.n187 9.0005
R8307 iovss.n226 iovss.n187 9.0005
R8308 iovss.n216 iovss.n187 9.0005
R8309 iovss.n228 iovss.n187 9.0005
R8310 iovss.n215 iovss.n187 9.0005
R8311 iovss.n230 iovss.n187 9.0005
R8312 iovss.n214 iovss.n187 9.0005
R8313 iovss.n232 iovss.n187 9.0005
R8314 iovss.n213 iovss.n187 9.0005
R8315 iovss.n234 iovss.n187 9.0005
R8316 iovss.n212 iovss.n187 9.0005
R8317 iovss.n236 iovss.n187 9.0005
R8318 iovss.n211 iovss.n187 9.0005
R8319 iovss.n237 iovss.n187 9.0005
R8320 iovss.n3429 iovss.n187 9.0005
R8321 iovss.n239 iovss.n187 9.0005
R8322 iovss.n210 iovss.n187 9.0005
R8323 iovss.n241 iovss.n187 9.0005
R8324 iovss.n209 iovss.n187 9.0005
R8325 iovss.n243 iovss.n187 9.0005
R8326 iovss.n208 iovss.n187 9.0005
R8327 iovss.n245 iovss.n187 9.0005
R8328 iovss.n207 iovss.n187 9.0005
R8329 iovss.n247 iovss.n187 9.0005
R8330 iovss.n206 iovss.n187 9.0005
R8331 iovss.n248 iovss.n187 9.0005
R8332 iovss.n205 iovss.n187 9.0005
R8333 iovss.n250 iovss.n187 9.0005
R8334 iovss.n204 iovss.n187 9.0005
R8335 iovss.n251 iovss.n187 9.0005
R8336 iovss.n253 iovss.n187 9.0005
R8337 iovss.n3427 iovss.n187 9.0005
R8338 iovss.n219 iovss.n182 9.0005
R8339 iovss.n222 iovss.n182 9.0005
R8340 iovss.n218 iovss.n182 9.0005
R8341 iovss.n224 iovss.n182 9.0005
R8342 iovss.n217 iovss.n182 9.0005
R8343 iovss.n226 iovss.n182 9.0005
R8344 iovss.n216 iovss.n182 9.0005
R8345 iovss.n228 iovss.n182 9.0005
R8346 iovss.n215 iovss.n182 9.0005
R8347 iovss.n230 iovss.n182 9.0005
R8348 iovss.n214 iovss.n182 9.0005
R8349 iovss.n232 iovss.n182 9.0005
R8350 iovss.n213 iovss.n182 9.0005
R8351 iovss.n234 iovss.n182 9.0005
R8352 iovss.n212 iovss.n182 9.0005
R8353 iovss.n236 iovss.n182 9.0005
R8354 iovss.n211 iovss.n182 9.0005
R8355 iovss.n237 iovss.n182 9.0005
R8356 iovss.n3429 iovss.n182 9.0005
R8357 iovss.n239 iovss.n182 9.0005
R8358 iovss.n210 iovss.n182 9.0005
R8359 iovss.n241 iovss.n182 9.0005
R8360 iovss.n209 iovss.n182 9.0005
R8361 iovss.n243 iovss.n182 9.0005
R8362 iovss.n208 iovss.n182 9.0005
R8363 iovss.n245 iovss.n182 9.0005
R8364 iovss.n207 iovss.n182 9.0005
R8365 iovss.n247 iovss.n182 9.0005
R8366 iovss.n206 iovss.n182 9.0005
R8367 iovss.n248 iovss.n182 9.0005
R8368 iovss.n205 iovss.n182 9.0005
R8369 iovss.n250 iovss.n182 9.0005
R8370 iovss.n204 iovss.n182 9.0005
R8371 iovss.n251 iovss.n182 9.0005
R8372 iovss.n253 iovss.n182 9.0005
R8373 iovss.n3427 iovss.n182 9.0005
R8374 iovss.n219 iovss.n188 9.0005
R8375 iovss.n222 iovss.n188 9.0005
R8376 iovss.n218 iovss.n188 9.0005
R8377 iovss.n224 iovss.n188 9.0005
R8378 iovss.n217 iovss.n188 9.0005
R8379 iovss.n226 iovss.n188 9.0005
R8380 iovss.n216 iovss.n188 9.0005
R8381 iovss.n228 iovss.n188 9.0005
R8382 iovss.n215 iovss.n188 9.0005
R8383 iovss.n230 iovss.n188 9.0005
R8384 iovss.n214 iovss.n188 9.0005
R8385 iovss.n232 iovss.n188 9.0005
R8386 iovss.n213 iovss.n188 9.0005
R8387 iovss.n234 iovss.n188 9.0005
R8388 iovss.n212 iovss.n188 9.0005
R8389 iovss.n236 iovss.n188 9.0005
R8390 iovss.n211 iovss.n188 9.0005
R8391 iovss.n237 iovss.n188 9.0005
R8392 iovss.n3429 iovss.n188 9.0005
R8393 iovss.n239 iovss.n188 9.0005
R8394 iovss.n210 iovss.n188 9.0005
R8395 iovss.n241 iovss.n188 9.0005
R8396 iovss.n209 iovss.n188 9.0005
R8397 iovss.n243 iovss.n188 9.0005
R8398 iovss.n208 iovss.n188 9.0005
R8399 iovss.n245 iovss.n188 9.0005
R8400 iovss.n207 iovss.n188 9.0005
R8401 iovss.n247 iovss.n188 9.0005
R8402 iovss.n206 iovss.n188 9.0005
R8403 iovss.n248 iovss.n188 9.0005
R8404 iovss.n205 iovss.n188 9.0005
R8405 iovss.n250 iovss.n188 9.0005
R8406 iovss.n204 iovss.n188 9.0005
R8407 iovss.n251 iovss.n188 9.0005
R8408 iovss.n253 iovss.n188 9.0005
R8409 iovss.n3427 iovss.n188 9.0005
R8410 iovss.n219 iovss.n181 9.0005
R8411 iovss.n222 iovss.n181 9.0005
R8412 iovss.n218 iovss.n181 9.0005
R8413 iovss.n224 iovss.n181 9.0005
R8414 iovss.n217 iovss.n181 9.0005
R8415 iovss.n226 iovss.n181 9.0005
R8416 iovss.n216 iovss.n181 9.0005
R8417 iovss.n228 iovss.n181 9.0005
R8418 iovss.n215 iovss.n181 9.0005
R8419 iovss.n230 iovss.n181 9.0005
R8420 iovss.n214 iovss.n181 9.0005
R8421 iovss.n232 iovss.n181 9.0005
R8422 iovss.n213 iovss.n181 9.0005
R8423 iovss.n234 iovss.n181 9.0005
R8424 iovss.n212 iovss.n181 9.0005
R8425 iovss.n236 iovss.n181 9.0005
R8426 iovss.n211 iovss.n181 9.0005
R8427 iovss.n237 iovss.n181 9.0005
R8428 iovss.n3429 iovss.n181 9.0005
R8429 iovss.n239 iovss.n181 9.0005
R8430 iovss.n210 iovss.n181 9.0005
R8431 iovss.n241 iovss.n181 9.0005
R8432 iovss.n209 iovss.n181 9.0005
R8433 iovss.n243 iovss.n181 9.0005
R8434 iovss.n208 iovss.n181 9.0005
R8435 iovss.n245 iovss.n181 9.0005
R8436 iovss.n207 iovss.n181 9.0005
R8437 iovss.n247 iovss.n181 9.0005
R8438 iovss.n206 iovss.n181 9.0005
R8439 iovss.n248 iovss.n181 9.0005
R8440 iovss.n205 iovss.n181 9.0005
R8441 iovss.n250 iovss.n181 9.0005
R8442 iovss.n204 iovss.n181 9.0005
R8443 iovss.n251 iovss.n181 9.0005
R8444 iovss.n253 iovss.n181 9.0005
R8445 iovss.n3427 iovss.n181 9.0005
R8446 iovss.n219 iovss.n189 9.0005
R8447 iovss.n222 iovss.n189 9.0005
R8448 iovss.n218 iovss.n189 9.0005
R8449 iovss.n224 iovss.n189 9.0005
R8450 iovss.n217 iovss.n189 9.0005
R8451 iovss.n226 iovss.n189 9.0005
R8452 iovss.n216 iovss.n189 9.0005
R8453 iovss.n228 iovss.n189 9.0005
R8454 iovss.n215 iovss.n189 9.0005
R8455 iovss.n230 iovss.n189 9.0005
R8456 iovss.n214 iovss.n189 9.0005
R8457 iovss.n232 iovss.n189 9.0005
R8458 iovss.n213 iovss.n189 9.0005
R8459 iovss.n234 iovss.n189 9.0005
R8460 iovss.n212 iovss.n189 9.0005
R8461 iovss.n236 iovss.n189 9.0005
R8462 iovss.n211 iovss.n189 9.0005
R8463 iovss.n237 iovss.n189 9.0005
R8464 iovss.n3429 iovss.n189 9.0005
R8465 iovss.n239 iovss.n189 9.0005
R8466 iovss.n210 iovss.n189 9.0005
R8467 iovss.n241 iovss.n189 9.0005
R8468 iovss.n209 iovss.n189 9.0005
R8469 iovss.n243 iovss.n189 9.0005
R8470 iovss.n208 iovss.n189 9.0005
R8471 iovss.n245 iovss.n189 9.0005
R8472 iovss.n207 iovss.n189 9.0005
R8473 iovss.n247 iovss.n189 9.0005
R8474 iovss.n206 iovss.n189 9.0005
R8475 iovss.n248 iovss.n189 9.0005
R8476 iovss.n205 iovss.n189 9.0005
R8477 iovss.n250 iovss.n189 9.0005
R8478 iovss.n204 iovss.n189 9.0005
R8479 iovss.n251 iovss.n189 9.0005
R8480 iovss.n253 iovss.n189 9.0005
R8481 iovss.n3427 iovss.n189 9.0005
R8482 iovss.n219 iovss.n180 9.0005
R8483 iovss.n222 iovss.n180 9.0005
R8484 iovss.n218 iovss.n180 9.0005
R8485 iovss.n224 iovss.n180 9.0005
R8486 iovss.n217 iovss.n180 9.0005
R8487 iovss.n226 iovss.n180 9.0005
R8488 iovss.n216 iovss.n180 9.0005
R8489 iovss.n228 iovss.n180 9.0005
R8490 iovss.n215 iovss.n180 9.0005
R8491 iovss.n230 iovss.n180 9.0005
R8492 iovss.n214 iovss.n180 9.0005
R8493 iovss.n232 iovss.n180 9.0005
R8494 iovss.n213 iovss.n180 9.0005
R8495 iovss.n234 iovss.n180 9.0005
R8496 iovss.n212 iovss.n180 9.0005
R8497 iovss.n236 iovss.n180 9.0005
R8498 iovss.n211 iovss.n180 9.0005
R8499 iovss.n237 iovss.n180 9.0005
R8500 iovss.n3429 iovss.n180 9.0005
R8501 iovss.n239 iovss.n180 9.0005
R8502 iovss.n210 iovss.n180 9.0005
R8503 iovss.n241 iovss.n180 9.0005
R8504 iovss.n209 iovss.n180 9.0005
R8505 iovss.n243 iovss.n180 9.0005
R8506 iovss.n208 iovss.n180 9.0005
R8507 iovss.n245 iovss.n180 9.0005
R8508 iovss.n207 iovss.n180 9.0005
R8509 iovss.n247 iovss.n180 9.0005
R8510 iovss.n206 iovss.n180 9.0005
R8511 iovss.n248 iovss.n180 9.0005
R8512 iovss.n205 iovss.n180 9.0005
R8513 iovss.n250 iovss.n180 9.0005
R8514 iovss.n204 iovss.n180 9.0005
R8515 iovss.n251 iovss.n180 9.0005
R8516 iovss.n253 iovss.n180 9.0005
R8517 iovss.n3427 iovss.n180 9.0005
R8518 iovss.n219 iovss.n190 9.0005
R8519 iovss.n222 iovss.n190 9.0005
R8520 iovss.n218 iovss.n190 9.0005
R8521 iovss.n224 iovss.n190 9.0005
R8522 iovss.n217 iovss.n190 9.0005
R8523 iovss.n226 iovss.n190 9.0005
R8524 iovss.n216 iovss.n190 9.0005
R8525 iovss.n228 iovss.n190 9.0005
R8526 iovss.n215 iovss.n190 9.0005
R8527 iovss.n230 iovss.n190 9.0005
R8528 iovss.n214 iovss.n190 9.0005
R8529 iovss.n232 iovss.n190 9.0005
R8530 iovss.n213 iovss.n190 9.0005
R8531 iovss.n234 iovss.n190 9.0005
R8532 iovss.n212 iovss.n190 9.0005
R8533 iovss.n236 iovss.n190 9.0005
R8534 iovss.n211 iovss.n190 9.0005
R8535 iovss.n237 iovss.n190 9.0005
R8536 iovss.n3429 iovss.n190 9.0005
R8537 iovss.n239 iovss.n190 9.0005
R8538 iovss.n210 iovss.n190 9.0005
R8539 iovss.n241 iovss.n190 9.0005
R8540 iovss.n209 iovss.n190 9.0005
R8541 iovss.n243 iovss.n190 9.0005
R8542 iovss.n208 iovss.n190 9.0005
R8543 iovss.n245 iovss.n190 9.0005
R8544 iovss.n207 iovss.n190 9.0005
R8545 iovss.n247 iovss.n190 9.0005
R8546 iovss.n206 iovss.n190 9.0005
R8547 iovss.n248 iovss.n190 9.0005
R8548 iovss.n205 iovss.n190 9.0005
R8549 iovss.n250 iovss.n190 9.0005
R8550 iovss.n204 iovss.n190 9.0005
R8551 iovss.n251 iovss.n190 9.0005
R8552 iovss.n253 iovss.n190 9.0005
R8553 iovss.n3427 iovss.n190 9.0005
R8554 iovss.n219 iovss.n179 9.0005
R8555 iovss.n222 iovss.n179 9.0005
R8556 iovss.n218 iovss.n179 9.0005
R8557 iovss.n224 iovss.n179 9.0005
R8558 iovss.n217 iovss.n179 9.0005
R8559 iovss.n226 iovss.n179 9.0005
R8560 iovss.n216 iovss.n179 9.0005
R8561 iovss.n228 iovss.n179 9.0005
R8562 iovss.n215 iovss.n179 9.0005
R8563 iovss.n230 iovss.n179 9.0005
R8564 iovss.n214 iovss.n179 9.0005
R8565 iovss.n232 iovss.n179 9.0005
R8566 iovss.n213 iovss.n179 9.0005
R8567 iovss.n234 iovss.n179 9.0005
R8568 iovss.n212 iovss.n179 9.0005
R8569 iovss.n236 iovss.n179 9.0005
R8570 iovss.n211 iovss.n179 9.0005
R8571 iovss.n237 iovss.n179 9.0005
R8572 iovss.n3429 iovss.n179 9.0005
R8573 iovss.n239 iovss.n179 9.0005
R8574 iovss.n210 iovss.n179 9.0005
R8575 iovss.n241 iovss.n179 9.0005
R8576 iovss.n209 iovss.n179 9.0005
R8577 iovss.n243 iovss.n179 9.0005
R8578 iovss.n208 iovss.n179 9.0005
R8579 iovss.n245 iovss.n179 9.0005
R8580 iovss.n207 iovss.n179 9.0005
R8581 iovss.n247 iovss.n179 9.0005
R8582 iovss.n206 iovss.n179 9.0005
R8583 iovss.n248 iovss.n179 9.0005
R8584 iovss.n205 iovss.n179 9.0005
R8585 iovss.n250 iovss.n179 9.0005
R8586 iovss.n204 iovss.n179 9.0005
R8587 iovss.n251 iovss.n179 9.0005
R8588 iovss.n253 iovss.n179 9.0005
R8589 iovss.n3427 iovss.n179 9.0005
R8590 iovss.n219 iovss.n191 9.0005
R8591 iovss.n222 iovss.n191 9.0005
R8592 iovss.n218 iovss.n191 9.0005
R8593 iovss.n224 iovss.n191 9.0005
R8594 iovss.n217 iovss.n191 9.0005
R8595 iovss.n226 iovss.n191 9.0005
R8596 iovss.n216 iovss.n191 9.0005
R8597 iovss.n228 iovss.n191 9.0005
R8598 iovss.n215 iovss.n191 9.0005
R8599 iovss.n230 iovss.n191 9.0005
R8600 iovss.n214 iovss.n191 9.0005
R8601 iovss.n232 iovss.n191 9.0005
R8602 iovss.n213 iovss.n191 9.0005
R8603 iovss.n234 iovss.n191 9.0005
R8604 iovss.n212 iovss.n191 9.0005
R8605 iovss.n236 iovss.n191 9.0005
R8606 iovss.n211 iovss.n191 9.0005
R8607 iovss.n237 iovss.n191 9.0005
R8608 iovss.n3429 iovss.n191 9.0005
R8609 iovss.n239 iovss.n191 9.0005
R8610 iovss.n210 iovss.n191 9.0005
R8611 iovss.n241 iovss.n191 9.0005
R8612 iovss.n209 iovss.n191 9.0005
R8613 iovss.n243 iovss.n191 9.0005
R8614 iovss.n208 iovss.n191 9.0005
R8615 iovss.n245 iovss.n191 9.0005
R8616 iovss.n207 iovss.n191 9.0005
R8617 iovss.n247 iovss.n191 9.0005
R8618 iovss.n206 iovss.n191 9.0005
R8619 iovss.n248 iovss.n191 9.0005
R8620 iovss.n205 iovss.n191 9.0005
R8621 iovss.n250 iovss.n191 9.0005
R8622 iovss.n204 iovss.n191 9.0005
R8623 iovss.n251 iovss.n191 9.0005
R8624 iovss.n253 iovss.n191 9.0005
R8625 iovss.n3427 iovss.n191 9.0005
R8626 iovss.n219 iovss.n178 9.0005
R8627 iovss.n222 iovss.n178 9.0005
R8628 iovss.n218 iovss.n178 9.0005
R8629 iovss.n224 iovss.n178 9.0005
R8630 iovss.n217 iovss.n178 9.0005
R8631 iovss.n226 iovss.n178 9.0005
R8632 iovss.n216 iovss.n178 9.0005
R8633 iovss.n228 iovss.n178 9.0005
R8634 iovss.n215 iovss.n178 9.0005
R8635 iovss.n230 iovss.n178 9.0005
R8636 iovss.n214 iovss.n178 9.0005
R8637 iovss.n232 iovss.n178 9.0005
R8638 iovss.n213 iovss.n178 9.0005
R8639 iovss.n234 iovss.n178 9.0005
R8640 iovss.n212 iovss.n178 9.0005
R8641 iovss.n236 iovss.n178 9.0005
R8642 iovss.n211 iovss.n178 9.0005
R8643 iovss.n237 iovss.n178 9.0005
R8644 iovss.n3429 iovss.n178 9.0005
R8645 iovss.n239 iovss.n178 9.0005
R8646 iovss.n210 iovss.n178 9.0005
R8647 iovss.n241 iovss.n178 9.0005
R8648 iovss.n209 iovss.n178 9.0005
R8649 iovss.n243 iovss.n178 9.0005
R8650 iovss.n208 iovss.n178 9.0005
R8651 iovss.n245 iovss.n178 9.0005
R8652 iovss.n207 iovss.n178 9.0005
R8653 iovss.n247 iovss.n178 9.0005
R8654 iovss.n206 iovss.n178 9.0005
R8655 iovss.n248 iovss.n178 9.0005
R8656 iovss.n205 iovss.n178 9.0005
R8657 iovss.n250 iovss.n178 9.0005
R8658 iovss.n204 iovss.n178 9.0005
R8659 iovss.n251 iovss.n178 9.0005
R8660 iovss.n253 iovss.n178 9.0005
R8661 iovss.n3427 iovss.n178 9.0005
R8662 iovss.n219 iovss.n192 9.0005
R8663 iovss.n222 iovss.n192 9.0005
R8664 iovss.n218 iovss.n192 9.0005
R8665 iovss.n224 iovss.n192 9.0005
R8666 iovss.n217 iovss.n192 9.0005
R8667 iovss.n226 iovss.n192 9.0005
R8668 iovss.n216 iovss.n192 9.0005
R8669 iovss.n228 iovss.n192 9.0005
R8670 iovss.n215 iovss.n192 9.0005
R8671 iovss.n230 iovss.n192 9.0005
R8672 iovss.n214 iovss.n192 9.0005
R8673 iovss.n232 iovss.n192 9.0005
R8674 iovss.n213 iovss.n192 9.0005
R8675 iovss.n234 iovss.n192 9.0005
R8676 iovss.n212 iovss.n192 9.0005
R8677 iovss.n236 iovss.n192 9.0005
R8678 iovss.n211 iovss.n192 9.0005
R8679 iovss.n237 iovss.n192 9.0005
R8680 iovss.n3429 iovss.n192 9.0005
R8681 iovss.n239 iovss.n192 9.0005
R8682 iovss.n210 iovss.n192 9.0005
R8683 iovss.n241 iovss.n192 9.0005
R8684 iovss.n209 iovss.n192 9.0005
R8685 iovss.n243 iovss.n192 9.0005
R8686 iovss.n208 iovss.n192 9.0005
R8687 iovss.n245 iovss.n192 9.0005
R8688 iovss.n207 iovss.n192 9.0005
R8689 iovss.n247 iovss.n192 9.0005
R8690 iovss.n206 iovss.n192 9.0005
R8691 iovss.n248 iovss.n192 9.0005
R8692 iovss.n205 iovss.n192 9.0005
R8693 iovss.n250 iovss.n192 9.0005
R8694 iovss.n204 iovss.n192 9.0005
R8695 iovss.n251 iovss.n192 9.0005
R8696 iovss.n253 iovss.n192 9.0005
R8697 iovss.n3427 iovss.n192 9.0005
R8698 iovss.n219 iovss.n177 9.0005
R8699 iovss.n222 iovss.n177 9.0005
R8700 iovss.n218 iovss.n177 9.0005
R8701 iovss.n224 iovss.n177 9.0005
R8702 iovss.n217 iovss.n177 9.0005
R8703 iovss.n226 iovss.n177 9.0005
R8704 iovss.n216 iovss.n177 9.0005
R8705 iovss.n228 iovss.n177 9.0005
R8706 iovss.n215 iovss.n177 9.0005
R8707 iovss.n230 iovss.n177 9.0005
R8708 iovss.n214 iovss.n177 9.0005
R8709 iovss.n232 iovss.n177 9.0005
R8710 iovss.n213 iovss.n177 9.0005
R8711 iovss.n234 iovss.n177 9.0005
R8712 iovss.n212 iovss.n177 9.0005
R8713 iovss.n236 iovss.n177 9.0005
R8714 iovss.n211 iovss.n177 9.0005
R8715 iovss.n237 iovss.n177 9.0005
R8716 iovss.n3429 iovss.n177 9.0005
R8717 iovss.n239 iovss.n177 9.0005
R8718 iovss.n210 iovss.n177 9.0005
R8719 iovss.n241 iovss.n177 9.0005
R8720 iovss.n209 iovss.n177 9.0005
R8721 iovss.n243 iovss.n177 9.0005
R8722 iovss.n208 iovss.n177 9.0005
R8723 iovss.n245 iovss.n177 9.0005
R8724 iovss.n207 iovss.n177 9.0005
R8725 iovss.n247 iovss.n177 9.0005
R8726 iovss.n206 iovss.n177 9.0005
R8727 iovss.n248 iovss.n177 9.0005
R8728 iovss.n205 iovss.n177 9.0005
R8729 iovss.n250 iovss.n177 9.0005
R8730 iovss.n204 iovss.n177 9.0005
R8731 iovss.n251 iovss.n177 9.0005
R8732 iovss.n253 iovss.n177 9.0005
R8733 iovss.n3427 iovss.n177 9.0005
R8734 iovss.n219 iovss.n193 9.0005
R8735 iovss.n222 iovss.n193 9.0005
R8736 iovss.n218 iovss.n193 9.0005
R8737 iovss.n224 iovss.n193 9.0005
R8738 iovss.n217 iovss.n193 9.0005
R8739 iovss.n226 iovss.n193 9.0005
R8740 iovss.n216 iovss.n193 9.0005
R8741 iovss.n228 iovss.n193 9.0005
R8742 iovss.n215 iovss.n193 9.0005
R8743 iovss.n230 iovss.n193 9.0005
R8744 iovss.n214 iovss.n193 9.0005
R8745 iovss.n232 iovss.n193 9.0005
R8746 iovss.n213 iovss.n193 9.0005
R8747 iovss.n234 iovss.n193 9.0005
R8748 iovss.n212 iovss.n193 9.0005
R8749 iovss.n236 iovss.n193 9.0005
R8750 iovss.n211 iovss.n193 9.0005
R8751 iovss.n237 iovss.n193 9.0005
R8752 iovss.n3429 iovss.n193 9.0005
R8753 iovss.n239 iovss.n193 9.0005
R8754 iovss.n210 iovss.n193 9.0005
R8755 iovss.n241 iovss.n193 9.0005
R8756 iovss.n209 iovss.n193 9.0005
R8757 iovss.n243 iovss.n193 9.0005
R8758 iovss.n208 iovss.n193 9.0005
R8759 iovss.n245 iovss.n193 9.0005
R8760 iovss.n207 iovss.n193 9.0005
R8761 iovss.n247 iovss.n193 9.0005
R8762 iovss.n206 iovss.n193 9.0005
R8763 iovss.n248 iovss.n193 9.0005
R8764 iovss.n205 iovss.n193 9.0005
R8765 iovss.n250 iovss.n193 9.0005
R8766 iovss.n204 iovss.n193 9.0005
R8767 iovss.n251 iovss.n193 9.0005
R8768 iovss.n253 iovss.n193 9.0005
R8769 iovss.n3427 iovss.n193 9.0005
R8770 iovss.n219 iovss.n176 9.0005
R8771 iovss.n222 iovss.n176 9.0005
R8772 iovss.n218 iovss.n176 9.0005
R8773 iovss.n224 iovss.n176 9.0005
R8774 iovss.n217 iovss.n176 9.0005
R8775 iovss.n226 iovss.n176 9.0005
R8776 iovss.n216 iovss.n176 9.0005
R8777 iovss.n228 iovss.n176 9.0005
R8778 iovss.n215 iovss.n176 9.0005
R8779 iovss.n230 iovss.n176 9.0005
R8780 iovss.n214 iovss.n176 9.0005
R8781 iovss.n232 iovss.n176 9.0005
R8782 iovss.n213 iovss.n176 9.0005
R8783 iovss.n234 iovss.n176 9.0005
R8784 iovss.n212 iovss.n176 9.0005
R8785 iovss.n236 iovss.n176 9.0005
R8786 iovss.n211 iovss.n176 9.0005
R8787 iovss.n237 iovss.n176 9.0005
R8788 iovss.n3429 iovss.n176 9.0005
R8789 iovss.n239 iovss.n176 9.0005
R8790 iovss.n210 iovss.n176 9.0005
R8791 iovss.n241 iovss.n176 9.0005
R8792 iovss.n209 iovss.n176 9.0005
R8793 iovss.n243 iovss.n176 9.0005
R8794 iovss.n208 iovss.n176 9.0005
R8795 iovss.n245 iovss.n176 9.0005
R8796 iovss.n207 iovss.n176 9.0005
R8797 iovss.n247 iovss.n176 9.0005
R8798 iovss.n206 iovss.n176 9.0005
R8799 iovss.n248 iovss.n176 9.0005
R8800 iovss.n205 iovss.n176 9.0005
R8801 iovss.n250 iovss.n176 9.0005
R8802 iovss.n204 iovss.n176 9.0005
R8803 iovss.n251 iovss.n176 9.0005
R8804 iovss.n253 iovss.n176 9.0005
R8805 iovss.n3427 iovss.n176 9.0005
R8806 iovss.n3428 iovss.n219 9.0005
R8807 iovss.n3428 iovss.n222 9.0005
R8808 iovss.n3428 iovss.n218 9.0005
R8809 iovss.n3428 iovss.n224 9.0005
R8810 iovss.n3428 iovss.n217 9.0005
R8811 iovss.n3428 iovss.n226 9.0005
R8812 iovss.n3428 iovss.n216 9.0005
R8813 iovss.n3428 iovss.n228 9.0005
R8814 iovss.n3428 iovss.n215 9.0005
R8815 iovss.n3428 iovss.n230 9.0005
R8816 iovss.n3428 iovss.n214 9.0005
R8817 iovss.n3428 iovss.n232 9.0005
R8818 iovss.n3428 iovss.n213 9.0005
R8819 iovss.n3428 iovss.n234 9.0005
R8820 iovss.n3428 iovss.n212 9.0005
R8821 iovss.n3428 iovss.n236 9.0005
R8822 iovss.n3428 iovss.n211 9.0005
R8823 iovss.n3428 iovss.n237 9.0005
R8824 iovss.n3429 iovss.n3428 9.0005
R8825 iovss.n3428 iovss.n239 9.0005
R8826 iovss.n3428 iovss.n210 9.0005
R8827 iovss.n3428 iovss.n241 9.0005
R8828 iovss.n3428 iovss.n209 9.0005
R8829 iovss.n3428 iovss.n243 9.0005
R8830 iovss.n3428 iovss.n208 9.0005
R8831 iovss.n3428 iovss.n245 9.0005
R8832 iovss.n3428 iovss.n207 9.0005
R8833 iovss.n3428 iovss.n247 9.0005
R8834 iovss.n3428 iovss.n206 9.0005
R8835 iovss.n3428 iovss.n248 9.0005
R8836 iovss.n3428 iovss.n205 9.0005
R8837 iovss.n3428 iovss.n250 9.0005
R8838 iovss.n3428 iovss.n204 9.0005
R8839 iovss.n3428 iovss.n251 9.0005
R8840 iovss.n3428 iovss.n203 9.0005
R8841 iovss.n3428 iovss.n253 9.0005
R8842 iovss.n3428 iovss.n3427 9.0005
R8843 iovss.n3394 iovss.n275 9.0005
R8844 iovss.n306 iovss.n275 9.0005
R8845 iovss.n301 iovss.n275 9.0005
R8846 iovss.n309 iovss.n275 9.0005
R8847 iovss.n299 iovss.n275 9.0005
R8848 iovss.n312 iovss.n275 9.0005
R8849 iovss.n297 iovss.n275 9.0005
R8850 iovss.n315 iovss.n275 9.0005
R8851 iovss.n295 iovss.n275 9.0005
R8852 iovss.n318 iovss.n275 9.0005
R8853 iovss.n293 iovss.n275 9.0005
R8854 iovss.n3390 iovss.n275 9.0005
R8855 iovss.n3392 iovss.n275 9.0005
R8856 iovss.n3391 iovss.n291 9.0005
R8857 iovss.n3391 iovss.n324 9.0005
R8858 iovss.n3391 iovss.n289 9.0005
R8859 iovss.n3391 iovss.n328 9.0005
R8860 iovss.n3391 iovss.n287 9.0005
R8861 iovss.n3391 iovss.n331 9.0005
R8862 iovss.n3391 iovss.n3390 9.0005
R8863 iovss.n3392 iovss.n3391 9.0005
R8864 iovss.n3394 iovss.n274 9.0005
R8865 iovss.n305 iovss.n274 9.0005
R8866 iovss.n302 iovss.n274 9.0005
R8867 iovss.n306 iovss.n274 9.0005
R8868 iovss.n301 iovss.n274 9.0005
R8869 iovss.n308 iovss.n274 9.0005
R8870 iovss.n300 iovss.n274 9.0005
R8871 iovss.n309 iovss.n274 9.0005
R8872 iovss.n299 iovss.n274 9.0005
R8873 iovss.n311 iovss.n274 9.0005
R8874 iovss.n298 iovss.n274 9.0005
R8875 iovss.n312 iovss.n274 9.0005
R8876 iovss.n297 iovss.n274 9.0005
R8877 iovss.n314 iovss.n274 9.0005
R8878 iovss.n296 iovss.n274 9.0005
R8879 iovss.n315 iovss.n274 9.0005
R8880 iovss.n295 iovss.n274 9.0005
R8881 iovss.n317 iovss.n274 9.0005
R8882 iovss.n294 iovss.n274 9.0005
R8883 iovss.n318 iovss.n274 9.0005
R8884 iovss.n293 iovss.n274 9.0005
R8885 iovss.n320 iovss.n274 9.0005
R8886 iovss.n292 iovss.n274 9.0005
R8887 iovss.n322 iovss.n274 9.0005
R8888 iovss.n291 iovss.n274 9.0005
R8889 iovss.n324 iovss.n274 9.0005
R8890 iovss.n290 iovss.n274 9.0005
R8891 iovss.n326 iovss.n274 9.0005
R8892 iovss.n289 iovss.n274 9.0005
R8893 iovss.n328 iovss.n274 9.0005
R8894 iovss.n288 iovss.n274 9.0005
R8895 iovss.n330 iovss.n274 9.0005
R8896 iovss.n287 iovss.n274 9.0005
R8897 iovss.n331 iovss.n274 9.0005
R8898 iovss.n3390 iovss.n274 9.0005
R8899 iovss.n3392 iovss.n274 9.0005
R8900 iovss.n3394 iovss.n277 9.0005
R8901 iovss.n305 iovss.n277 9.0005
R8902 iovss.n302 iovss.n277 9.0005
R8903 iovss.n306 iovss.n277 9.0005
R8904 iovss.n301 iovss.n277 9.0005
R8905 iovss.n308 iovss.n277 9.0005
R8906 iovss.n300 iovss.n277 9.0005
R8907 iovss.n309 iovss.n277 9.0005
R8908 iovss.n299 iovss.n277 9.0005
R8909 iovss.n311 iovss.n277 9.0005
R8910 iovss.n298 iovss.n277 9.0005
R8911 iovss.n312 iovss.n277 9.0005
R8912 iovss.n297 iovss.n277 9.0005
R8913 iovss.n314 iovss.n277 9.0005
R8914 iovss.n296 iovss.n277 9.0005
R8915 iovss.n315 iovss.n277 9.0005
R8916 iovss.n295 iovss.n277 9.0005
R8917 iovss.n317 iovss.n277 9.0005
R8918 iovss.n294 iovss.n277 9.0005
R8919 iovss.n318 iovss.n277 9.0005
R8920 iovss.n293 iovss.n277 9.0005
R8921 iovss.n320 iovss.n277 9.0005
R8922 iovss.n292 iovss.n277 9.0005
R8923 iovss.n322 iovss.n277 9.0005
R8924 iovss.n291 iovss.n277 9.0005
R8925 iovss.n324 iovss.n277 9.0005
R8926 iovss.n290 iovss.n277 9.0005
R8927 iovss.n326 iovss.n277 9.0005
R8928 iovss.n289 iovss.n277 9.0005
R8929 iovss.n328 iovss.n277 9.0005
R8930 iovss.n288 iovss.n277 9.0005
R8931 iovss.n330 iovss.n277 9.0005
R8932 iovss.n287 iovss.n277 9.0005
R8933 iovss.n331 iovss.n277 9.0005
R8934 iovss.n3390 iovss.n277 9.0005
R8935 iovss.n3392 iovss.n277 9.0005
R8936 iovss.n3394 iovss.n273 9.0005
R8937 iovss.n305 iovss.n273 9.0005
R8938 iovss.n302 iovss.n273 9.0005
R8939 iovss.n306 iovss.n273 9.0005
R8940 iovss.n301 iovss.n273 9.0005
R8941 iovss.n308 iovss.n273 9.0005
R8942 iovss.n300 iovss.n273 9.0005
R8943 iovss.n309 iovss.n273 9.0005
R8944 iovss.n299 iovss.n273 9.0005
R8945 iovss.n311 iovss.n273 9.0005
R8946 iovss.n298 iovss.n273 9.0005
R8947 iovss.n312 iovss.n273 9.0005
R8948 iovss.n297 iovss.n273 9.0005
R8949 iovss.n314 iovss.n273 9.0005
R8950 iovss.n296 iovss.n273 9.0005
R8951 iovss.n315 iovss.n273 9.0005
R8952 iovss.n295 iovss.n273 9.0005
R8953 iovss.n317 iovss.n273 9.0005
R8954 iovss.n294 iovss.n273 9.0005
R8955 iovss.n318 iovss.n273 9.0005
R8956 iovss.n293 iovss.n273 9.0005
R8957 iovss.n320 iovss.n273 9.0005
R8958 iovss.n292 iovss.n273 9.0005
R8959 iovss.n322 iovss.n273 9.0005
R8960 iovss.n291 iovss.n273 9.0005
R8961 iovss.n324 iovss.n273 9.0005
R8962 iovss.n290 iovss.n273 9.0005
R8963 iovss.n326 iovss.n273 9.0005
R8964 iovss.n289 iovss.n273 9.0005
R8965 iovss.n328 iovss.n273 9.0005
R8966 iovss.n288 iovss.n273 9.0005
R8967 iovss.n330 iovss.n273 9.0005
R8968 iovss.n287 iovss.n273 9.0005
R8969 iovss.n331 iovss.n273 9.0005
R8970 iovss.n3390 iovss.n273 9.0005
R8971 iovss.n3392 iovss.n273 9.0005
R8972 iovss.n3394 iovss.n278 9.0005
R8973 iovss.n305 iovss.n278 9.0005
R8974 iovss.n302 iovss.n278 9.0005
R8975 iovss.n306 iovss.n278 9.0005
R8976 iovss.n301 iovss.n278 9.0005
R8977 iovss.n308 iovss.n278 9.0005
R8978 iovss.n300 iovss.n278 9.0005
R8979 iovss.n309 iovss.n278 9.0005
R8980 iovss.n299 iovss.n278 9.0005
R8981 iovss.n311 iovss.n278 9.0005
R8982 iovss.n298 iovss.n278 9.0005
R8983 iovss.n312 iovss.n278 9.0005
R8984 iovss.n297 iovss.n278 9.0005
R8985 iovss.n314 iovss.n278 9.0005
R8986 iovss.n296 iovss.n278 9.0005
R8987 iovss.n315 iovss.n278 9.0005
R8988 iovss.n295 iovss.n278 9.0005
R8989 iovss.n317 iovss.n278 9.0005
R8990 iovss.n294 iovss.n278 9.0005
R8991 iovss.n318 iovss.n278 9.0005
R8992 iovss.n293 iovss.n278 9.0005
R8993 iovss.n320 iovss.n278 9.0005
R8994 iovss.n292 iovss.n278 9.0005
R8995 iovss.n322 iovss.n278 9.0005
R8996 iovss.n291 iovss.n278 9.0005
R8997 iovss.n324 iovss.n278 9.0005
R8998 iovss.n290 iovss.n278 9.0005
R8999 iovss.n326 iovss.n278 9.0005
R9000 iovss.n289 iovss.n278 9.0005
R9001 iovss.n328 iovss.n278 9.0005
R9002 iovss.n288 iovss.n278 9.0005
R9003 iovss.n330 iovss.n278 9.0005
R9004 iovss.n287 iovss.n278 9.0005
R9005 iovss.n331 iovss.n278 9.0005
R9006 iovss.n3390 iovss.n278 9.0005
R9007 iovss.n3392 iovss.n278 9.0005
R9008 iovss.n3394 iovss.n272 9.0005
R9009 iovss.n305 iovss.n272 9.0005
R9010 iovss.n302 iovss.n272 9.0005
R9011 iovss.n306 iovss.n272 9.0005
R9012 iovss.n301 iovss.n272 9.0005
R9013 iovss.n308 iovss.n272 9.0005
R9014 iovss.n300 iovss.n272 9.0005
R9015 iovss.n309 iovss.n272 9.0005
R9016 iovss.n299 iovss.n272 9.0005
R9017 iovss.n311 iovss.n272 9.0005
R9018 iovss.n298 iovss.n272 9.0005
R9019 iovss.n312 iovss.n272 9.0005
R9020 iovss.n297 iovss.n272 9.0005
R9021 iovss.n314 iovss.n272 9.0005
R9022 iovss.n296 iovss.n272 9.0005
R9023 iovss.n315 iovss.n272 9.0005
R9024 iovss.n295 iovss.n272 9.0005
R9025 iovss.n317 iovss.n272 9.0005
R9026 iovss.n294 iovss.n272 9.0005
R9027 iovss.n318 iovss.n272 9.0005
R9028 iovss.n293 iovss.n272 9.0005
R9029 iovss.n320 iovss.n272 9.0005
R9030 iovss.n292 iovss.n272 9.0005
R9031 iovss.n322 iovss.n272 9.0005
R9032 iovss.n291 iovss.n272 9.0005
R9033 iovss.n324 iovss.n272 9.0005
R9034 iovss.n290 iovss.n272 9.0005
R9035 iovss.n326 iovss.n272 9.0005
R9036 iovss.n289 iovss.n272 9.0005
R9037 iovss.n328 iovss.n272 9.0005
R9038 iovss.n288 iovss.n272 9.0005
R9039 iovss.n330 iovss.n272 9.0005
R9040 iovss.n287 iovss.n272 9.0005
R9041 iovss.n331 iovss.n272 9.0005
R9042 iovss.n3390 iovss.n272 9.0005
R9043 iovss.n3392 iovss.n272 9.0005
R9044 iovss.n3394 iovss.n279 9.0005
R9045 iovss.n305 iovss.n279 9.0005
R9046 iovss.n302 iovss.n279 9.0005
R9047 iovss.n306 iovss.n279 9.0005
R9048 iovss.n301 iovss.n279 9.0005
R9049 iovss.n308 iovss.n279 9.0005
R9050 iovss.n300 iovss.n279 9.0005
R9051 iovss.n309 iovss.n279 9.0005
R9052 iovss.n299 iovss.n279 9.0005
R9053 iovss.n311 iovss.n279 9.0005
R9054 iovss.n298 iovss.n279 9.0005
R9055 iovss.n312 iovss.n279 9.0005
R9056 iovss.n297 iovss.n279 9.0005
R9057 iovss.n314 iovss.n279 9.0005
R9058 iovss.n296 iovss.n279 9.0005
R9059 iovss.n315 iovss.n279 9.0005
R9060 iovss.n295 iovss.n279 9.0005
R9061 iovss.n317 iovss.n279 9.0005
R9062 iovss.n294 iovss.n279 9.0005
R9063 iovss.n318 iovss.n279 9.0005
R9064 iovss.n293 iovss.n279 9.0005
R9065 iovss.n320 iovss.n279 9.0005
R9066 iovss.n292 iovss.n279 9.0005
R9067 iovss.n322 iovss.n279 9.0005
R9068 iovss.n291 iovss.n279 9.0005
R9069 iovss.n324 iovss.n279 9.0005
R9070 iovss.n290 iovss.n279 9.0005
R9071 iovss.n326 iovss.n279 9.0005
R9072 iovss.n289 iovss.n279 9.0005
R9073 iovss.n328 iovss.n279 9.0005
R9074 iovss.n288 iovss.n279 9.0005
R9075 iovss.n330 iovss.n279 9.0005
R9076 iovss.n287 iovss.n279 9.0005
R9077 iovss.n331 iovss.n279 9.0005
R9078 iovss.n3390 iovss.n279 9.0005
R9079 iovss.n3392 iovss.n279 9.0005
R9080 iovss.n3394 iovss.n271 9.0005
R9081 iovss.n305 iovss.n271 9.0005
R9082 iovss.n302 iovss.n271 9.0005
R9083 iovss.n306 iovss.n271 9.0005
R9084 iovss.n301 iovss.n271 9.0005
R9085 iovss.n308 iovss.n271 9.0005
R9086 iovss.n300 iovss.n271 9.0005
R9087 iovss.n309 iovss.n271 9.0005
R9088 iovss.n299 iovss.n271 9.0005
R9089 iovss.n311 iovss.n271 9.0005
R9090 iovss.n298 iovss.n271 9.0005
R9091 iovss.n312 iovss.n271 9.0005
R9092 iovss.n297 iovss.n271 9.0005
R9093 iovss.n314 iovss.n271 9.0005
R9094 iovss.n296 iovss.n271 9.0005
R9095 iovss.n315 iovss.n271 9.0005
R9096 iovss.n295 iovss.n271 9.0005
R9097 iovss.n317 iovss.n271 9.0005
R9098 iovss.n294 iovss.n271 9.0005
R9099 iovss.n318 iovss.n271 9.0005
R9100 iovss.n293 iovss.n271 9.0005
R9101 iovss.n320 iovss.n271 9.0005
R9102 iovss.n292 iovss.n271 9.0005
R9103 iovss.n322 iovss.n271 9.0005
R9104 iovss.n291 iovss.n271 9.0005
R9105 iovss.n324 iovss.n271 9.0005
R9106 iovss.n290 iovss.n271 9.0005
R9107 iovss.n326 iovss.n271 9.0005
R9108 iovss.n289 iovss.n271 9.0005
R9109 iovss.n328 iovss.n271 9.0005
R9110 iovss.n288 iovss.n271 9.0005
R9111 iovss.n330 iovss.n271 9.0005
R9112 iovss.n287 iovss.n271 9.0005
R9113 iovss.n331 iovss.n271 9.0005
R9114 iovss.n3390 iovss.n271 9.0005
R9115 iovss.n3392 iovss.n271 9.0005
R9116 iovss.n3394 iovss.n280 9.0005
R9117 iovss.n305 iovss.n280 9.0005
R9118 iovss.n302 iovss.n280 9.0005
R9119 iovss.n306 iovss.n280 9.0005
R9120 iovss.n301 iovss.n280 9.0005
R9121 iovss.n308 iovss.n280 9.0005
R9122 iovss.n300 iovss.n280 9.0005
R9123 iovss.n309 iovss.n280 9.0005
R9124 iovss.n299 iovss.n280 9.0005
R9125 iovss.n311 iovss.n280 9.0005
R9126 iovss.n298 iovss.n280 9.0005
R9127 iovss.n312 iovss.n280 9.0005
R9128 iovss.n297 iovss.n280 9.0005
R9129 iovss.n314 iovss.n280 9.0005
R9130 iovss.n296 iovss.n280 9.0005
R9131 iovss.n315 iovss.n280 9.0005
R9132 iovss.n295 iovss.n280 9.0005
R9133 iovss.n317 iovss.n280 9.0005
R9134 iovss.n294 iovss.n280 9.0005
R9135 iovss.n318 iovss.n280 9.0005
R9136 iovss.n293 iovss.n280 9.0005
R9137 iovss.n320 iovss.n280 9.0005
R9138 iovss.n292 iovss.n280 9.0005
R9139 iovss.n322 iovss.n280 9.0005
R9140 iovss.n291 iovss.n280 9.0005
R9141 iovss.n324 iovss.n280 9.0005
R9142 iovss.n290 iovss.n280 9.0005
R9143 iovss.n326 iovss.n280 9.0005
R9144 iovss.n289 iovss.n280 9.0005
R9145 iovss.n328 iovss.n280 9.0005
R9146 iovss.n288 iovss.n280 9.0005
R9147 iovss.n330 iovss.n280 9.0005
R9148 iovss.n287 iovss.n280 9.0005
R9149 iovss.n331 iovss.n280 9.0005
R9150 iovss.n3390 iovss.n280 9.0005
R9151 iovss.n3392 iovss.n280 9.0005
R9152 iovss.n3394 iovss.n270 9.0005
R9153 iovss.n305 iovss.n270 9.0005
R9154 iovss.n302 iovss.n270 9.0005
R9155 iovss.n306 iovss.n270 9.0005
R9156 iovss.n301 iovss.n270 9.0005
R9157 iovss.n308 iovss.n270 9.0005
R9158 iovss.n300 iovss.n270 9.0005
R9159 iovss.n309 iovss.n270 9.0005
R9160 iovss.n299 iovss.n270 9.0005
R9161 iovss.n311 iovss.n270 9.0005
R9162 iovss.n298 iovss.n270 9.0005
R9163 iovss.n312 iovss.n270 9.0005
R9164 iovss.n297 iovss.n270 9.0005
R9165 iovss.n314 iovss.n270 9.0005
R9166 iovss.n296 iovss.n270 9.0005
R9167 iovss.n315 iovss.n270 9.0005
R9168 iovss.n295 iovss.n270 9.0005
R9169 iovss.n317 iovss.n270 9.0005
R9170 iovss.n294 iovss.n270 9.0005
R9171 iovss.n318 iovss.n270 9.0005
R9172 iovss.n293 iovss.n270 9.0005
R9173 iovss.n320 iovss.n270 9.0005
R9174 iovss.n292 iovss.n270 9.0005
R9175 iovss.n322 iovss.n270 9.0005
R9176 iovss.n291 iovss.n270 9.0005
R9177 iovss.n324 iovss.n270 9.0005
R9178 iovss.n290 iovss.n270 9.0005
R9179 iovss.n326 iovss.n270 9.0005
R9180 iovss.n289 iovss.n270 9.0005
R9181 iovss.n328 iovss.n270 9.0005
R9182 iovss.n288 iovss.n270 9.0005
R9183 iovss.n330 iovss.n270 9.0005
R9184 iovss.n287 iovss.n270 9.0005
R9185 iovss.n331 iovss.n270 9.0005
R9186 iovss.n3390 iovss.n270 9.0005
R9187 iovss.n3392 iovss.n270 9.0005
R9188 iovss.n3394 iovss.n281 9.0005
R9189 iovss.n305 iovss.n281 9.0005
R9190 iovss.n302 iovss.n281 9.0005
R9191 iovss.n306 iovss.n281 9.0005
R9192 iovss.n301 iovss.n281 9.0005
R9193 iovss.n308 iovss.n281 9.0005
R9194 iovss.n300 iovss.n281 9.0005
R9195 iovss.n309 iovss.n281 9.0005
R9196 iovss.n299 iovss.n281 9.0005
R9197 iovss.n311 iovss.n281 9.0005
R9198 iovss.n298 iovss.n281 9.0005
R9199 iovss.n312 iovss.n281 9.0005
R9200 iovss.n297 iovss.n281 9.0005
R9201 iovss.n314 iovss.n281 9.0005
R9202 iovss.n296 iovss.n281 9.0005
R9203 iovss.n315 iovss.n281 9.0005
R9204 iovss.n295 iovss.n281 9.0005
R9205 iovss.n317 iovss.n281 9.0005
R9206 iovss.n294 iovss.n281 9.0005
R9207 iovss.n318 iovss.n281 9.0005
R9208 iovss.n293 iovss.n281 9.0005
R9209 iovss.n320 iovss.n281 9.0005
R9210 iovss.n292 iovss.n281 9.0005
R9211 iovss.n322 iovss.n281 9.0005
R9212 iovss.n291 iovss.n281 9.0005
R9213 iovss.n324 iovss.n281 9.0005
R9214 iovss.n290 iovss.n281 9.0005
R9215 iovss.n326 iovss.n281 9.0005
R9216 iovss.n289 iovss.n281 9.0005
R9217 iovss.n328 iovss.n281 9.0005
R9218 iovss.n288 iovss.n281 9.0005
R9219 iovss.n330 iovss.n281 9.0005
R9220 iovss.n287 iovss.n281 9.0005
R9221 iovss.n331 iovss.n281 9.0005
R9222 iovss.n3390 iovss.n281 9.0005
R9223 iovss.n3392 iovss.n281 9.0005
R9224 iovss.n3394 iovss.n269 9.0005
R9225 iovss.n305 iovss.n269 9.0005
R9226 iovss.n302 iovss.n269 9.0005
R9227 iovss.n306 iovss.n269 9.0005
R9228 iovss.n301 iovss.n269 9.0005
R9229 iovss.n308 iovss.n269 9.0005
R9230 iovss.n300 iovss.n269 9.0005
R9231 iovss.n309 iovss.n269 9.0005
R9232 iovss.n299 iovss.n269 9.0005
R9233 iovss.n311 iovss.n269 9.0005
R9234 iovss.n298 iovss.n269 9.0005
R9235 iovss.n312 iovss.n269 9.0005
R9236 iovss.n297 iovss.n269 9.0005
R9237 iovss.n314 iovss.n269 9.0005
R9238 iovss.n296 iovss.n269 9.0005
R9239 iovss.n315 iovss.n269 9.0005
R9240 iovss.n295 iovss.n269 9.0005
R9241 iovss.n317 iovss.n269 9.0005
R9242 iovss.n294 iovss.n269 9.0005
R9243 iovss.n318 iovss.n269 9.0005
R9244 iovss.n293 iovss.n269 9.0005
R9245 iovss.n320 iovss.n269 9.0005
R9246 iovss.n292 iovss.n269 9.0005
R9247 iovss.n322 iovss.n269 9.0005
R9248 iovss.n291 iovss.n269 9.0005
R9249 iovss.n324 iovss.n269 9.0005
R9250 iovss.n290 iovss.n269 9.0005
R9251 iovss.n326 iovss.n269 9.0005
R9252 iovss.n289 iovss.n269 9.0005
R9253 iovss.n328 iovss.n269 9.0005
R9254 iovss.n288 iovss.n269 9.0005
R9255 iovss.n330 iovss.n269 9.0005
R9256 iovss.n287 iovss.n269 9.0005
R9257 iovss.n331 iovss.n269 9.0005
R9258 iovss.n3390 iovss.n269 9.0005
R9259 iovss.n3392 iovss.n269 9.0005
R9260 iovss.n3394 iovss.n282 9.0005
R9261 iovss.n305 iovss.n282 9.0005
R9262 iovss.n302 iovss.n282 9.0005
R9263 iovss.n306 iovss.n282 9.0005
R9264 iovss.n301 iovss.n282 9.0005
R9265 iovss.n308 iovss.n282 9.0005
R9266 iovss.n300 iovss.n282 9.0005
R9267 iovss.n309 iovss.n282 9.0005
R9268 iovss.n299 iovss.n282 9.0005
R9269 iovss.n311 iovss.n282 9.0005
R9270 iovss.n298 iovss.n282 9.0005
R9271 iovss.n312 iovss.n282 9.0005
R9272 iovss.n297 iovss.n282 9.0005
R9273 iovss.n314 iovss.n282 9.0005
R9274 iovss.n296 iovss.n282 9.0005
R9275 iovss.n315 iovss.n282 9.0005
R9276 iovss.n295 iovss.n282 9.0005
R9277 iovss.n317 iovss.n282 9.0005
R9278 iovss.n294 iovss.n282 9.0005
R9279 iovss.n318 iovss.n282 9.0005
R9280 iovss.n293 iovss.n282 9.0005
R9281 iovss.n320 iovss.n282 9.0005
R9282 iovss.n292 iovss.n282 9.0005
R9283 iovss.n322 iovss.n282 9.0005
R9284 iovss.n291 iovss.n282 9.0005
R9285 iovss.n324 iovss.n282 9.0005
R9286 iovss.n290 iovss.n282 9.0005
R9287 iovss.n326 iovss.n282 9.0005
R9288 iovss.n289 iovss.n282 9.0005
R9289 iovss.n328 iovss.n282 9.0005
R9290 iovss.n288 iovss.n282 9.0005
R9291 iovss.n330 iovss.n282 9.0005
R9292 iovss.n287 iovss.n282 9.0005
R9293 iovss.n331 iovss.n282 9.0005
R9294 iovss.n3390 iovss.n282 9.0005
R9295 iovss.n3392 iovss.n282 9.0005
R9296 iovss.n3394 iovss.n268 9.0005
R9297 iovss.n305 iovss.n268 9.0005
R9298 iovss.n302 iovss.n268 9.0005
R9299 iovss.n306 iovss.n268 9.0005
R9300 iovss.n301 iovss.n268 9.0005
R9301 iovss.n308 iovss.n268 9.0005
R9302 iovss.n300 iovss.n268 9.0005
R9303 iovss.n309 iovss.n268 9.0005
R9304 iovss.n299 iovss.n268 9.0005
R9305 iovss.n311 iovss.n268 9.0005
R9306 iovss.n298 iovss.n268 9.0005
R9307 iovss.n312 iovss.n268 9.0005
R9308 iovss.n297 iovss.n268 9.0005
R9309 iovss.n314 iovss.n268 9.0005
R9310 iovss.n296 iovss.n268 9.0005
R9311 iovss.n315 iovss.n268 9.0005
R9312 iovss.n295 iovss.n268 9.0005
R9313 iovss.n317 iovss.n268 9.0005
R9314 iovss.n294 iovss.n268 9.0005
R9315 iovss.n318 iovss.n268 9.0005
R9316 iovss.n293 iovss.n268 9.0005
R9317 iovss.n320 iovss.n268 9.0005
R9318 iovss.n292 iovss.n268 9.0005
R9319 iovss.n322 iovss.n268 9.0005
R9320 iovss.n291 iovss.n268 9.0005
R9321 iovss.n324 iovss.n268 9.0005
R9322 iovss.n290 iovss.n268 9.0005
R9323 iovss.n326 iovss.n268 9.0005
R9324 iovss.n289 iovss.n268 9.0005
R9325 iovss.n328 iovss.n268 9.0005
R9326 iovss.n288 iovss.n268 9.0005
R9327 iovss.n330 iovss.n268 9.0005
R9328 iovss.n287 iovss.n268 9.0005
R9329 iovss.n331 iovss.n268 9.0005
R9330 iovss.n3390 iovss.n268 9.0005
R9331 iovss.n3392 iovss.n268 9.0005
R9332 iovss.n3394 iovss.n283 9.0005
R9333 iovss.n305 iovss.n283 9.0005
R9334 iovss.n302 iovss.n283 9.0005
R9335 iovss.n306 iovss.n283 9.0005
R9336 iovss.n301 iovss.n283 9.0005
R9337 iovss.n308 iovss.n283 9.0005
R9338 iovss.n300 iovss.n283 9.0005
R9339 iovss.n309 iovss.n283 9.0005
R9340 iovss.n299 iovss.n283 9.0005
R9341 iovss.n311 iovss.n283 9.0005
R9342 iovss.n298 iovss.n283 9.0005
R9343 iovss.n312 iovss.n283 9.0005
R9344 iovss.n297 iovss.n283 9.0005
R9345 iovss.n314 iovss.n283 9.0005
R9346 iovss.n296 iovss.n283 9.0005
R9347 iovss.n315 iovss.n283 9.0005
R9348 iovss.n295 iovss.n283 9.0005
R9349 iovss.n317 iovss.n283 9.0005
R9350 iovss.n294 iovss.n283 9.0005
R9351 iovss.n318 iovss.n283 9.0005
R9352 iovss.n293 iovss.n283 9.0005
R9353 iovss.n320 iovss.n283 9.0005
R9354 iovss.n292 iovss.n283 9.0005
R9355 iovss.n322 iovss.n283 9.0005
R9356 iovss.n291 iovss.n283 9.0005
R9357 iovss.n324 iovss.n283 9.0005
R9358 iovss.n290 iovss.n283 9.0005
R9359 iovss.n326 iovss.n283 9.0005
R9360 iovss.n289 iovss.n283 9.0005
R9361 iovss.n328 iovss.n283 9.0005
R9362 iovss.n288 iovss.n283 9.0005
R9363 iovss.n330 iovss.n283 9.0005
R9364 iovss.n287 iovss.n283 9.0005
R9365 iovss.n331 iovss.n283 9.0005
R9366 iovss.n3390 iovss.n283 9.0005
R9367 iovss.n3392 iovss.n283 9.0005
R9368 iovss.n3394 iovss.n267 9.0005
R9369 iovss.n305 iovss.n267 9.0005
R9370 iovss.n302 iovss.n267 9.0005
R9371 iovss.n306 iovss.n267 9.0005
R9372 iovss.n301 iovss.n267 9.0005
R9373 iovss.n308 iovss.n267 9.0005
R9374 iovss.n300 iovss.n267 9.0005
R9375 iovss.n309 iovss.n267 9.0005
R9376 iovss.n299 iovss.n267 9.0005
R9377 iovss.n311 iovss.n267 9.0005
R9378 iovss.n298 iovss.n267 9.0005
R9379 iovss.n312 iovss.n267 9.0005
R9380 iovss.n297 iovss.n267 9.0005
R9381 iovss.n314 iovss.n267 9.0005
R9382 iovss.n296 iovss.n267 9.0005
R9383 iovss.n315 iovss.n267 9.0005
R9384 iovss.n295 iovss.n267 9.0005
R9385 iovss.n317 iovss.n267 9.0005
R9386 iovss.n294 iovss.n267 9.0005
R9387 iovss.n318 iovss.n267 9.0005
R9388 iovss.n293 iovss.n267 9.0005
R9389 iovss.n320 iovss.n267 9.0005
R9390 iovss.n292 iovss.n267 9.0005
R9391 iovss.n322 iovss.n267 9.0005
R9392 iovss.n291 iovss.n267 9.0005
R9393 iovss.n324 iovss.n267 9.0005
R9394 iovss.n290 iovss.n267 9.0005
R9395 iovss.n326 iovss.n267 9.0005
R9396 iovss.n289 iovss.n267 9.0005
R9397 iovss.n328 iovss.n267 9.0005
R9398 iovss.n288 iovss.n267 9.0005
R9399 iovss.n330 iovss.n267 9.0005
R9400 iovss.n287 iovss.n267 9.0005
R9401 iovss.n331 iovss.n267 9.0005
R9402 iovss.n3390 iovss.n267 9.0005
R9403 iovss.n3392 iovss.n267 9.0005
R9404 iovss.n3394 iovss.n284 9.0005
R9405 iovss.n305 iovss.n284 9.0005
R9406 iovss.n302 iovss.n284 9.0005
R9407 iovss.n306 iovss.n284 9.0005
R9408 iovss.n301 iovss.n284 9.0005
R9409 iovss.n308 iovss.n284 9.0005
R9410 iovss.n300 iovss.n284 9.0005
R9411 iovss.n309 iovss.n284 9.0005
R9412 iovss.n299 iovss.n284 9.0005
R9413 iovss.n311 iovss.n284 9.0005
R9414 iovss.n298 iovss.n284 9.0005
R9415 iovss.n312 iovss.n284 9.0005
R9416 iovss.n297 iovss.n284 9.0005
R9417 iovss.n314 iovss.n284 9.0005
R9418 iovss.n296 iovss.n284 9.0005
R9419 iovss.n315 iovss.n284 9.0005
R9420 iovss.n295 iovss.n284 9.0005
R9421 iovss.n317 iovss.n284 9.0005
R9422 iovss.n294 iovss.n284 9.0005
R9423 iovss.n318 iovss.n284 9.0005
R9424 iovss.n293 iovss.n284 9.0005
R9425 iovss.n320 iovss.n284 9.0005
R9426 iovss.n292 iovss.n284 9.0005
R9427 iovss.n322 iovss.n284 9.0005
R9428 iovss.n291 iovss.n284 9.0005
R9429 iovss.n324 iovss.n284 9.0005
R9430 iovss.n290 iovss.n284 9.0005
R9431 iovss.n326 iovss.n284 9.0005
R9432 iovss.n289 iovss.n284 9.0005
R9433 iovss.n328 iovss.n284 9.0005
R9434 iovss.n288 iovss.n284 9.0005
R9435 iovss.n330 iovss.n284 9.0005
R9436 iovss.n287 iovss.n284 9.0005
R9437 iovss.n331 iovss.n284 9.0005
R9438 iovss.n3390 iovss.n284 9.0005
R9439 iovss.n3392 iovss.n284 9.0005
R9440 iovss.n3394 iovss.n266 9.0005
R9441 iovss.n305 iovss.n266 9.0005
R9442 iovss.n302 iovss.n266 9.0005
R9443 iovss.n306 iovss.n266 9.0005
R9444 iovss.n301 iovss.n266 9.0005
R9445 iovss.n308 iovss.n266 9.0005
R9446 iovss.n300 iovss.n266 9.0005
R9447 iovss.n309 iovss.n266 9.0005
R9448 iovss.n299 iovss.n266 9.0005
R9449 iovss.n311 iovss.n266 9.0005
R9450 iovss.n298 iovss.n266 9.0005
R9451 iovss.n312 iovss.n266 9.0005
R9452 iovss.n297 iovss.n266 9.0005
R9453 iovss.n314 iovss.n266 9.0005
R9454 iovss.n296 iovss.n266 9.0005
R9455 iovss.n315 iovss.n266 9.0005
R9456 iovss.n295 iovss.n266 9.0005
R9457 iovss.n317 iovss.n266 9.0005
R9458 iovss.n294 iovss.n266 9.0005
R9459 iovss.n318 iovss.n266 9.0005
R9460 iovss.n293 iovss.n266 9.0005
R9461 iovss.n320 iovss.n266 9.0005
R9462 iovss.n292 iovss.n266 9.0005
R9463 iovss.n322 iovss.n266 9.0005
R9464 iovss.n291 iovss.n266 9.0005
R9465 iovss.n324 iovss.n266 9.0005
R9466 iovss.n290 iovss.n266 9.0005
R9467 iovss.n326 iovss.n266 9.0005
R9468 iovss.n289 iovss.n266 9.0005
R9469 iovss.n328 iovss.n266 9.0005
R9470 iovss.n288 iovss.n266 9.0005
R9471 iovss.n330 iovss.n266 9.0005
R9472 iovss.n287 iovss.n266 9.0005
R9473 iovss.n331 iovss.n266 9.0005
R9474 iovss.n3390 iovss.n266 9.0005
R9475 iovss.n3392 iovss.n266 9.0005
R9476 iovss.n3394 iovss.n3393 9.0005
R9477 iovss.n3393 iovss.n305 9.0005
R9478 iovss.n3393 iovss.n302 9.0005
R9479 iovss.n3393 iovss.n306 9.0005
R9480 iovss.n3393 iovss.n301 9.0005
R9481 iovss.n3393 iovss.n308 9.0005
R9482 iovss.n3393 iovss.n300 9.0005
R9483 iovss.n3393 iovss.n309 9.0005
R9484 iovss.n3393 iovss.n299 9.0005
R9485 iovss.n3393 iovss.n311 9.0005
R9486 iovss.n3393 iovss.n298 9.0005
R9487 iovss.n3393 iovss.n312 9.0005
R9488 iovss.n3393 iovss.n297 9.0005
R9489 iovss.n3393 iovss.n314 9.0005
R9490 iovss.n3393 iovss.n296 9.0005
R9491 iovss.n3393 iovss.n315 9.0005
R9492 iovss.n3393 iovss.n295 9.0005
R9493 iovss.n3393 iovss.n317 9.0005
R9494 iovss.n3393 iovss.n294 9.0005
R9495 iovss.n3393 iovss.n318 9.0005
R9496 iovss.n3393 iovss.n293 9.0005
R9497 iovss.n3393 iovss.n320 9.0005
R9498 iovss.n3393 iovss.n292 9.0005
R9499 iovss.n3393 iovss.n322 9.0005
R9500 iovss.n3393 iovss.n291 9.0005
R9501 iovss.n3393 iovss.n324 9.0005
R9502 iovss.n3393 iovss.n290 9.0005
R9503 iovss.n3393 iovss.n326 9.0005
R9504 iovss.n3393 iovss.n289 9.0005
R9505 iovss.n3393 iovss.n328 9.0005
R9506 iovss.n3393 iovss.n288 9.0005
R9507 iovss.n3393 iovss.n330 9.0005
R9508 iovss.n3393 iovss.n287 9.0005
R9509 iovss.n3393 iovss.n331 9.0005
R9510 iovss.n3393 iovss.n3392 9.0005
R9511 iovss.n672 iovss.n632 9.0005
R9512 iovss.n719 iovss.n632 9.0005
R9513 iovss.n661 iovss.n632 9.0005
R9514 iovss.n724 iovss.n632 9.0005
R9515 iovss.n659 iovss.n632 9.0005
R9516 iovss.n729 iovss.n632 9.0005
R9517 iovss.n657 iovss.n632 9.0005
R9518 iovss.n3246 iovss.n632 9.0005
R9519 iovss.n3249 iovss.n632 9.0005
R9520 iovss.n671 iovss.n646 9.0005
R9521 iovss.n678 iovss.n646 9.0005
R9522 iovss.n669 iovss.n646 9.0005
R9523 iovss.n683 iovss.n646 9.0005
R9524 iovss.n667 iovss.n646 9.0005
R9525 iovss.n688 iovss.n646 9.0005
R9526 iovss.n665 iovss.n646 9.0005
R9527 iovss.n710 iovss.n646 9.0005
R9528 iovss.n3251 iovss.n646 9.0005
R9529 iovss.n714 iovss.n646 9.0005
R9530 iovss.n3246 iovss.n646 9.0005
R9531 iovss.n3249 iovss.n646 9.0005
R9532 iovss.n672 iovss.n644 9.0005
R9533 iovss.n676 iovss.n644 9.0005
R9534 iovss.n671 iovss.n644 9.0005
R9535 iovss.n678 iovss.n644 9.0005
R9536 iovss.n670 iovss.n644 9.0005
R9537 iovss.n681 iovss.n644 9.0005
R9538 iovss.n669 iovss.n644 9.0005
R9539 iovss.n683 iovss.n644 9.0005
R9540 iovss.n668 iovss.n644 9.0005
R9541 iovss.n686 iovss.n644 9.0005
R9542 iovss.n667 iovss.n644 9.0005
R9543 iovss.n688 iovss.n644 9.0005
R9544 iovss.n666 iovss.n644 9.0005
R9545 iovss.n691 iovss.n644 9.0005
R9546 iovss.n665 iovss.n644 9.0005
R9547 iovss.n710 iovss.n644 9.0005
R9548 iovss.n664 iovss.n644 9.0005
R9549 iovss.n712 iovss.n644 9.0005
R9550 iovss.n3251 iovss.n644 9.0005
R9551 iovss.n714 iovss.n644 9.0005
R9552 iovss.n663 iovss.n644 9.0005
R9553 iovss.n717 iovss.n644 9.0005
R9554 iovss.n662 iovss.n644 9.0005
R9555 iovss.n719 iovss.n644 9.0005
R9556 iovss.n661 iovss.n644 9.0005
R9557 iovss.n722 iovss.n644 9.0005
R9558 iovss.n660 iovss.n644 9.0005
R9559 iovss.n724 iovss.n644 9.0005
R9560 iovss.n659 iovss.n644 9.0005
R9561 iovss.n727 iovss.n644 9.0005
R9562 iovss.n658 iovss.n644 9.0005
R9563 iovss.n729 iovss.n644 9.0005
R9564 iovss.n657 iovss.n644 9.0005
R9565 iovss.n731 iovss.n644 9.0005
R9566 iovss.n3246 iovss.n644 9.0005
R9567 iovss.n3249 iovss.n644 9.0005
R9568 iovss.n672 iovss.n647 9.0005
R9569 iovss.n676 iovss.n647 9.0005
R9570 iovss.n671 iovss.n647 9.0005
R9571 iovss.n678 iovss.n647 9.0005
R9572 iovss.n670 iovss.n647 9.0005
R9573 iovss.n681 iovss.n647 9.0005
R9574 iovss.n669 iovss.n647 9.0005
R9575 iovss.n683 iovss.n647 9.0005
R9576 iovss.n668 iovss.n647 9.0005
R9577 iovss.n686 iovss.n647 9.0005
R9578 iovss.n667 iovss.n647 9.0005
R9579 iovss.n688 iovss.n647 9.0005
R9580 iovss.n666 iovss.n647 9.0005
R9581 iovss.n691 iovss.n647 9.0005
R9582 iovss.n665 iovss.n647 9.0005
R9583 iovss.n710 iovss.n647 9.0005
R9584 iovss.n664 iovss.n647 9.0005
R9585 iovss.n712 iovss.n647 9.0005
R9586 iovss.n3251 iovss.n647 9.0005
R9587 iovss.n714 iovss.n647 9.0005
R9588 iovss.n663 iovss.n647 9.0005
R9589 iovss.n717 iovss.n647 9.0005
R9590 iovss.n662 iovss.n647 9.0005
R9591 iovss.n719 iovss.n647 9.0005
R9592 iovss.n661 iovss.n647 9.0005
R9593 iovss.n722 iovss.n647 9.0005
R9594 iovss.n660 iovss.n647 9.0005
R9595 iovss.n724 iovss.n647 9.0005
R9596 iovss.n659 iovss.n647 9.0005
R9597 iovss.n727 iovss.n647 9.0005
R9598 iovss.n658 iovss.n647 9.0005
R9599 iovss.n729 iovss.n647 9.0005
R9600 iovss.n657 iovss.n647 9.0005
R9601 iovss.n731 iovss.n647 9.0005
R9602 iovss.n3246 iovss.n647 9.0005
R9603 iovss.n3249 iovss.n647 9.0005
R9604 iovss.n672 iovss.n643 9.0005
R9605 iovss.n676 iovss.n643 9.0005
R9606 iovss.n671 iovss.n643 9.0005
R9607 iovss.n678 iovss.n643 9.0005
R9608 iovss.n670 iovss.n643 9.0005
R9609 iovss.n681 iovss.n643 9.0005
R9610 iovss.n669 iovss.n643 9.0005
R9611 iovss.n683 iovss.n643 9.0005
R9612 iovss.n668 iovss.n643 9.0005
R9613 iovss.n686 iovss.n643 9.0005
R9614 iovss.n667 iovss.n643 9.0005
R9615 iovss.n688 iovss.n643 9.0005
R9616 iovss.n666 iovss.n643 9.0005
R9617 iovss.n691 iovss.n643 9.0005
R9618 iovss.n665 iovss.n643 9.0005
R9619 iovss.n710 iovss.n643 9.0005
R9620 iovss.n664 iovss.n643 9.0005
R9621 iovss.n712 iovss.n643 9.0005
R9622 iovss.n3251 iovss.n643 9.0005
R9623 iovss.n714 iovss.n643 9.0005
R9624 iovss.n663 iovss.n643 9.0005
R9625 iovss.n717 iovss.n643 9.0005
R9626 iovss.n662 iovss.n643 9.0005
R9627 iovss.n719 iovss.n643 9.0005
R9628 iovss.n661 iovss.n643 9.0005
R9629 iovss.n722 iovss.n643 9.0005
R9630 iovss.n660 iovss.n643 9.0005
R9631 iovss.n724 iovss.n643 9.0005
R9632 iovss.n659 iovss.n643 9.0005
R9633 iovss.n727 iovss.n643 9.0005
R9634 iovss.n658 iovss.n643 9.0005
R9635 iovss.n729 iovss.n643 9.0005
R9636 iovss.n657 iovss.n643 9.0005
R9637 iovss.n731 iovss.n643 9.0005
R9638 iovss.n3246 iovss.n643 9.0005
R9639 iovss.n3249 iovss.n643 9.0005
R9640 iovss.n672 iovss.n648 9.0005
R9641 iovss.n676 iovss.n648 9.0005
R9642 iovss.n671 iovss.n648 9.0005
R9643 iovss.n678 iovss.n648 9.0005
R9644 iovss.n670 iovss.n648 9.0005
R9645 iovss.n681 iovss.n648 9.0005
R9646 iovss.n669 iovss.n648 9.0005
R9647 iovss.n683 iovss.n648 9.0005
R9648 iovss.n668 iovss.n648 9.0005
R9649 iovss.n686 iovss.n648 9.0005
R9650 iovss.n667 iovss.n648 9.0005
R9651 iovss.n688 iovss.n648 9.0005
R9652 iovss.n666 iovss.n648 9.0005
R9653 iovss.n691 iovss.n648 9.0005
R9654 iovss.n665 iovss.n648 9.0005
R9655 iovss.n710 iovss.n648 9.0005
R9656 iovss.n664 iovss.n648 9.0005
R9657 iovss.n712 iovss.n648 9.0005
R9658 iovss.n3251 iovss.n648 9.0005
R9659 iovss.n714 iovss.n648 9.0005
R9660 iovss.n663 iovss.n648 9.0005
R9661 iovss.n717 iovss.n648 9.0005
R9662 iovss.n662 iovss.n648 9.0005
R9663 iovss.n719 iovss.n648 9.0005
R9664 iovss.n661 iovss.n648 9.0005
R9665 iovss.n722 iovss.n648 9.0005
R9666 iovss.n660 iovss.n648 9.0005
R9667 iovss.n724 iovss.n648 9.0005
R9668 iovss.n659 iovss.n648 9.0005
R9669 iovss.n727 iovss.n648 9.0005
R9670 iovss.n658 iovss.n648 9.0005
R9671 iovss.n729 iovss.n648 9.0005
R9672 iovss.n657 iovss.n648 9.0005
R9673 iovss.n731 iovss.n648 9.0005
R9674 iovss.n3246 iovss.n648 9.0005
R9675 iovss.n3249 iovss.n648 9.0005
R9676 iovss.n672 iovss.n642 9.0005
R9677 iovss.n676 iovss.n642 9.0005
R9678 iovss.n671 iovss.n642 9.0005
R9679 iovss.n678 iovss.n642 9.0005
R9680 iovss.n670 iovss.n642 9.0005
R9681 iovss.n681 iovss.n642 9.0005
R9682 iovss.n669 iovss.n642 9.0005
R9683 iovss.n683 iovss.n642 9.0005
R9684 iovss.n668 iovss.n642 9.0005
R9685 iovss.n686 iovss.n642 9.0005
R9686 iovss.n667 iovss.n642 9.0005
R9687 iovss.n688 iovss.n642 9.0005
R9688 iovss.n666 iovss.n642 9.0005
R9689 iovss.n691 iovss.n642 9.0005
R9690 iovss.n665 iovss.n642 9.0005
R9691 iovss.n710 iovss.n642 9.0005
R9692 iovss.n664 iovss.n642 9.0005
R9693 iovss.n712 iovss.n642 9.0005
R9694 iovss.n3251 iovss.n642 9.0005
R9695 iovss.n714 iovss.n642 9.0005
R9696 iovss.n663 iovss.n642 9.0005
R9697 iovss.n717 iovss.n642 9.0005
R9698 iovss.n662 iovss.n642 9.0005
R9699 iovss.n719 iovss.n642 9.0005
R9700 iovss.n661 iovss.n642 9.0005
R9701 iovss.n722 iovss.n642 9.0005
R9702 iovss.n660 iovss.n642 9.0005
R9703 iovss.n724 iovss.n642 9.0005
R9704 iovss.n659 iovss.n642 9.0005
R9705 iovss.n727 iovss.n642 9.0005
R9706 iovss.n658 iovss.n642 9.0005
R9707 iovss.n729 iovss.n642 9.0005
R9708 iovss.n657 iovss.n642 9.0005
R9709 iovss.n731 iovss.n642 9.0005
R9710 iovss.n3246 iovss.n642 9.0005
R9711 iovss.n3249 iovss.n642 9.0005
R9712 iovss.n672 iovss.n649 9.0005
R9713 iovss.n676 iovss.n649 9.0005
R9714 iovss.n671 iovss.n649 9.0005
R9715 iovss.n678 iovss.n649 9.0005
R9716 iovss.n670 iovss.n649 9.0005
R9717 iovss.n681 iovss.n649 9.0005
R9718 iovss.n669 iovss.n649 9.0005
R9719 iovss.n683 iovss.n649 9.0005
R9720 iovss.n668 iovss.n649 9.0005
R9721 iovss.n686 iovss.n649 9.0005
R9722 iovss.n667 iovss.n649 9.0005
R9723 iovss.n688 iovss.n649 9.0005
R9724 iovss.n666 iovss.n649 9.0005
R9725 iovss.n691 iovss.n649 9.0005
R9726 iovss.n665 iovss.n649 9.0005
R9727 iovss.n710 iovss.n649 9.0005
R9728 iovss.n664 iovss.n649 9.0005
R9729 iovss.n712 iovss.n649 9.0005
R9730 iovss.n3251 iovss.n649 9.0005
R9731 iovss.n714 iovss.n649 9.0005
R9732 iovss.n663 iovss.n649 9.0005
R9733 iovss.n717 iovss.n649 9.0005
R9734 iovss.n662 iovss.n649 9.0005
R9735 iovss.n719 iovss.n649 9.0005
R9736 iovss.n661 iovss.n649 9.0005
R9737 iovss.n722 iovss.n649 9.0005
R9738 iovss.n660 iovss.n649 9.0005
R9739 iovss.n724 iovss.n649 9.0005
R9740 iovss.n659 iovss.n649 9.0005
R9741 iovss.n727 iovss.n649 9.0005
R9742 iovss.n658 iovss.n649 9.0005
R9743 iovss.n729 iovss.n649 9.0005
R9744 iovss.n657 iovss.n649 9.0005
R9745 iovss.n731 iovss.n649 9.0005
R9746 iovss.n3246 iovss.n649 9.0005
R9747 iovss.n3249 iovss.n649 9.0005
R9748 iovss.n672 iovss.n641 9.0005
R9749 iovss.n676 iovss.n641 9.0005
R9750 iovss.n671 iovss.n641 9.0005
R9751 iovss.n678 iovss.n641 9.0005
R9752 iovss.n670 iovss.n641 9.0005
R9753 iovss.n681 iovss.n641 9.0005
R9754 iovss.n669 iovss.n641 9.0005
R9755 iovss.n683 iovss.n641 9.0005
R9756 iovss.n668 iovss.n641 9.0005
R9757 iovss.n686 iovss.n641 9.0005
R9758 iovss.n667 iovss.n641 9.0005
R9759 iovss.n688 iovss.n641 9.0005
R9760 iovss.n666 iovss.n641 9.0005
R9761 iovss.n691 iovss.n641 9.0005
R9762 iovss.n665 iovss.n641 9.0005
R9763 iovss.n710 iovss.n641 9.0005
R9764 iovss.n664 iovss.n641 9.0005
R9765 iovss.n712 iovss.n641 9.0005
R9766 iovss.n3251 iovss.n641 9.0005
R9767 iovss.n714 iovss.n641 9.0005
R9768 iovss.n663 iovss.n641 9.0005
R9769 iovss.n717 iovss.n641 9.0005
R9770 iovss.n662 iovss.n641 9.0005
R9771 iovss.n719 iovss.n641 9.0005
R9772 iovss.n661 iovss.n641 9.0005
R9773 iovss.n722 iovss.n641 9.0005
R9774 iovss.n660 iovss.n641 9.0005
R9775 iovss.n724 iovss.n641 9.0005
R9776 iovss.n659 iovss.n641 9.0005
R9777 iovss.n727 iovss.n641 9.0005
R9778 iovss.n658 iovss.n641 9.0005
R9779 iovss.n729 iovss.n641 9.0005
R9780 iovss.n657 iovss.n641 9.0005
R9781 iovss.n731 iovss.n641 9.0005
R9782 iovss.n3246 iovss.n641 9.0005
R9783 iovss.n3249 iovss.n641 9.0005
R9784 iovss.n672 iovss.n650 9.0005
R9785 iovss.n676 iovss.n650 9.0005
R9786 iovss.n671 iovss.n650 9.0005
R9787 iovss.n678 iovss.n650 9.0005
R9788 iovss.n670 iovss.n650 9.0005
R9789 iovss.n681 iovss.n650 9.0005
R9790 iovss.n669 iovss.n650 9.0005
R9791 iovss.n683 iovss.n650 9.0005
R9792 iovss.n668 iovss.n650 9.0005
R9793 iovss.n686 iovss.n650 9.0005
R9794 iovss.n667 iovss.n650 9.0005
R9795 iovss.n688 iovss.n650 9.0005
R9796 iovss.n666 iovss.n650 9.0005
R9797 iovss.n691 iovss.n650 9.0005
R9798 iovss.n665 iovss.n650 9.0005
R9799 iovss.n710 iovss.n650 9.0005
R9800 iovss.n664 iovss.n650 9.0005
R9801 iovss.n712 iovss.n650 9.0005
R9802 iovss.n3251 iovss.n650 9.0005
R9803 iovss.n714 iovss.n650 9.0005
R9804 iovss.n663 iovss.n650 9.0005
R9805 iovss.n717 iovss.n650 9.0005
R9806 iovss.n662 iovss.n650 9.0005
R9807 iovss.n719 iovss.n650 9.0005
R9808 iovss.n661 iovss.n650 9.0005
R9809 iovss.n722 iovss.n650 9.0005
R9810 iovss.n660 iovss.n650 9.0005
R9811 iovss.n724 iovss.n650 9.0005
R9812 iovss.n659 iovss.n650 9.0005
R9813 iovss.n727 iovss.n650 9.0005
R9814 iovss.n658 iovss.n650 9.0005
R9815 iovss.n729 iovss.n650 9.0005
R9816 iovss.n657 iovss.n650 9.0005
R9817 iovss.n731 iovss.n650 9.0005
R9818 iovss.n3246 iovss.n650 9.0005
R9819 iovss.n3249 iovss.n650 9.0005
R9820 iovss.n672 iovss.n640 9.0005
R9821 iovss.n676 iovss.n640 9.0005
R9822 iovss.n671 iovss.n640 9.0005
R9823 iovss.n678 iovss.n640 9.0005
R9824 iovss.n670 iovss.n640 9.0005
R9825 iovss.n681 iovss.n640 9.0005
R9826 iovss.n669 iovss.n640 9.0005
R9827 iovss.n683 iovss.n640 9.0005
R9828 iovss.n668 iovss.n640 9.0005
R9829 iovss.n686 iovss.n640 9.0005
R9830 iovss.n667 iovss.n640 9.0005
R9831 iovss.n688 iovss.n640 9.0005
R9832 iovss.n666 iovss.n640 9.0005
R9833 iovss.n691 iovss.n640 9.0005
R9834 iovss.n665 iovss.n640 9.0005
R9835 iovss.n710 iovss.n640 9.0005
R9836 iovss.n664 iovss.n640 9.0005
R9837 iovss.n712 iovss.n640 9.0005
R9838 iovss.n3251 iovss.n640 9.0005
R9839 iovss.n714 iovss.n640 9.0005
R9840 iovss.n663 iovss.n640 9.0005
R9841 iovss.n717 iovss.n640 9.0005
R9842 iovss.n662 iovss.n640 9.0005
R9843 iovss.n719 iovss.n640 9.0005
R9844 iovss.n661 iovss.n640 9.0005
R9845 iovss.n722 iovss.n640 9.0005
R9846 iovss.n660 iovss.n640 9.0005
R9847 iovss.n724 iovss.n640 9.0005
R9848 iovss.n659 iovss.n640 9.0005
R9849 iovss.n727 iovss.n640 9.0005
R9850 iovss.n658 iovss.n640 9.0005
R9851 iovss.n729 iovss.n640 9.0005
R9852 iovss.n657 iovss.n640 9.0005
R9853 iovss.n731 iovss.n640 9.0005
R9854 iovss.n3246 iovss.n640 9.0005
R9855 iovss.n3249 iovss.n640 9.0005
R9856 iovss.n672 iovss.n651 9.0005
R9857 iovss.n676 iovss.n651 9.0005
R9858 iovss.n671 iovss.n651 9.0005
R9859 iovss.n678 iovss.n651 9.0005
R9860 iovss.n670 iovss.n651 9.0005
R9861 iovss.n681 iovss.n651 9.0005
R9862 iovss.n669 iovss.n651 9.0005
R9863 iovss.n683 iovss.n651 9.0005
R9864 iovss.n668 iovss.n651 9.0005
R9865 iovss.n686 iovss.n651 9.0005
R9866 iovss.n667 iovss.n651 9.0005
R9867 iovss.n688 iovss.n651 9.0005
R9868 iovss.n666 iovss.n651 9.0005
R9869 iovss.n691 iovss.n651 9.0005
R9870 iovss.n665 iovss.n651 9.0005
R9871 iovss.n710 iovss.n651 9.0005
R9872 iovss.n664 iovss.n651 9.0005
R9873 iovss.n712 iovss.n651 9.0005
R9874 iovss.n3251 iovss.n651 9.0005
R9875 iovss.n714 iovss.n651 9.0005
R9876 iovss.n663 iovss.n651 9.0005
R9877 iovss.n717 iovss.n651 9.0005
R9878 iovss.n662 iovss.n651 9.0005
R9879 iovss.n719 iovss.n651 9.0005
R9880 iovss.n661 iovss.n651 9.0005
R9881 iovss.n722 iovss.n651 9.0005
R9882 iovss.n660 iovss.n651 9.0005
R9883 iovss.n724 iovss.n651 9.0005
R9884 iovss.n659 iovss.n651 9.0005
R9885 iovss.n727 iovss.n651 9.0005
R9886 iovss.n658 iovss.n651 9.0005
R9887 iovss.n729 iovss.n651 9.0005
R9888 iovss.n657 iovss.n651 9.0005
R9889 iovss.n731 iovss.n651 9.0005
R9890 iovss.n3246 iovss.n651 9.0005
R9891 iovss.n3249 iovss.n651 9.0005
R9892 iovss.n672 iovss.n639 9.0005
R9893 iovss.n676 iovss.n639 9.0005
R9894 iovss.n671 iovss.n639 9.0005
R9895 iovss.n678 iovss.n639 9.0005
R9896 iovss.n670 iovss.n639 9.0005
R9897 iovss.n681 iovss.n639 9.0005
R9898 iovss.n669 iovss.n639 9.0005
R9899 iovss.n683 iovss.n639 9.0005
R9900 iovss.n668 iovss.n639 9.0005
R9901 iovss.n686 iovss.n639 9.0005
R9902 iovss.n667 iovss.n639 9.0005
R9903 iovss.n688 iovss.n639 9.0005
R9904 iovss.n666 iovss.n639 9.0005
R9905 iovss.n691 iovss.n639 9.0005
R9906 iovss.n665 iovss.n639 9.0005
R9907 iovss.n710 iovss.n639 9.0005
R9908 iovss.n664 iovss.n639 9.0005
R9909 iovss.n712 iovss.n639 9.0005
R9910 iovss.n3251 iovss.n639 9.0005
R9911 iovss.n714 iovss.n639 9.0005
R9912 iovss.n663 iovss.n639 9.0005
R9913 iovss.n717 iovss.n639 9.0005
R9914 iovss.n662 iovss.n639 9.0005
R9915 iovss.n719 iovss.n639 9.0005
R9916 iovss.n661 iovss.n639 9.0005
R9917 iovss.n722 iovss.n639 9.0005
R9918 iovss.n660 iovss.n639 9.0005
R9919 iovss.n724 iovss.n639 9.0005
R9920 iovss.n659 iovss.n639 9.0005
R9921 iovss.n727 iovss.n639 9.0005
R9922 iovss.n658 iovss.n639 9.0005
R9923 iovss.n729 iovss.n639 9.0005
R9924 iovss.n657 iovss.n639 9.0005
R9925 iovss.n731 iovss.n639 9.0005
R9926 iovss.n3246 iovss.n639 9.0005
R9927 iovss.n3249 iovss.n639 9.0005
R9928 iovss.n672 iovss.n652 9.0005
R9929 iovss.n676 iovss.n652 9.0005
R9930 iovss.n671 iovss.n652 9.0005
R9931 iovss.n678 iovss.n652 9.0005
R9932 iovss.n670 iovss.n652 9.0005
R9933 iovss.n681 iovss.n652 9.0005
R9934 iovss.n669 iovss.n652 9.0005
R9935 iovss.n683 iovss.n652 9.0005
R9936 iovss.n668 iovss.n652 9.0005
R9937 iovss.n686 iovss.n652 9.0005
R9938 iovss.n667 iovss.n652 9.0005
R9939 iovss.n688 iovss.n652 9.0005
R9940 iovss.n666 iovss.n652 9.0005
R9941 iovss.n691 iovss.n652 9.0005
R9942 iovss.n665 iovss.n652 9.0005
R9943 iovss.n710 iovss.n652 9.0005
R9944 iovss.n664 iovss.n652 9.0005
R9945 iovss.n712 iovss.n652 9.0005
R9946 iovss.n3251 iovss.n652 9.0005
R9947 iovss.n714 iovss.n652 9.0005
R9948 iovss.n663 iovss.n652 9.0005
R9949 iovss.n717 iovss.n652 9.0005
R9950 iovss.n662 iovss.n652 9.0005
R9951 iovss.n719 iovss.n652 9.0005
R9952 iovss.n661 iovss.n652 9.0005
R9953 iovss.n722 iovss.n652 9.0005
R9954 iovss.n660 iovss.n652 9.0005
R9955 iovss.n724 iovss.n652 9.0005
R9956 iovss.n659 iovss.n652 9.0005
R9957 iovss.n727 iovss.n652 9.0005
R9958 iovss.n658 iovss.n652 9.0005
R9959 iovss.n729 iovss.n652 9.0005
R9960 iovss.n657 iovss.n652 9.0005
R9961 iovss.n731 iovss.n652 9.0005
R9962 iovss.n3246 iovss.n652 9.0005
R9963 iovss.n3249 iovss.n652 9.0005
R9964 iovss.n672 iovss.n638 9.0005
R9965 iovss.n676 iovss.n638 9.0005
R9966 iovss.n671 iovss.n638 9.0005
R9967 iovss.n678 iovss.n638 9.0005
R9968 iovss.n670 iovss.n638 9.0005
R9969 iovss.n681 iovss.n638 9.0005
R9970 iovss.n669 iovss.n638 9.0005
R9971 iovss.n683 iovss.n638 9.0005
R9972 iovss.n668 iovss.n638 9.0005
R9973 iovss.n686 iovss.n638 9.0005
R9974 iovss.n667 iovss.n638 9.0005
R9975 iovss.n688 iovss.n638 9.0005
R9976 iovss.n666 iovss.n638 9.0005
R9977 iovss.n691 iovss.n638 9.0005
R9978 iovss.n665 iovss.n638 9.0005
R9979 iovss.n710 iovss.n638 9.0005
R9980 iovss.n664 iovss.n638 9.0005
R9981 iovss.n712 iovss.n638 9.0005
R9982 iovss.n3251 iovss.n638 9.0005
R9983 iovss.n714 iovss.n638 9.0005
R9984 iovss.n663 iovss.n638 9.0005
R9985 iovss.n717 iovss.n638 9.0005
R9986 iovss.n662 iovss.n638 9.0005
R9987 iovss.n719 iovss.n638 9.0005
R9988 iovss.n661 iovss.n638 9.0005
R9989 iovss.n722 iovss.n638 9.0005
R9990 iovss.n660 iovss.n638 9.0005
R9991 iovss.n724 iovss.n638 9.0005
R9992 iovss.n659 iovss.n638 9.0005
R9993 iovss.n727 iovss.n638 9.0005
R9994 iovss.n658 iovss.n638 9.0005
R9995 iovss.n729 iovss.n638 9.0005
R9996 iovss.n657 iovss.n638 9.0005
R9997 iovss.n731 iovss.n638 9.0005
R9998 iovss.n3246 iovss.n638 9.0005
R9999 iovss.n3249 iovss.n638 9.0005
R10000 iovss.n672 iovss.n653 9.0005
R10001 iovss.n676 iovss.n653 9.0005
R10002 iovss.n671 iovss.n653 9.0005
R10003 iovss.n678 iovss.n653 9.0005
R10004 iovss.n670 iovss.n653 9.0005
R10005 iovss.n681 iovss.n653 9.0005
R10006 iovss.n669 iovss.n653 9.0005
R10007 iovss.n683 iovss.n653 9.0005
R10008 iovss.n668 iovss.n653 9.0005
R10009 iovss.n686 iovss.n653 9.0005
R10010 iovss.n667 iovss.n653 9.0005
R10011 iovss.n688 iovss.n653 9.0005
R10012 iovss.n666 iovss.n653 9.0005
R10013 iovss.n691 iovss.n653 9.0005
R10014 iovss.n665 iovss.n653 9.0005
R10015 iovss.n710 iovss.n653 9.0005
R10016 iovss.n664 iovss.n653 9.0005
R10017 iovss.n712 iovss.n653 9.0005
R10018 iovss.n3251 iovss.n653 9.0005
R10019 iovss.n714 iovss.n653 9.0005
R10020 iovss.n663 iovss.n653 9.0005
R10021 iovss.n717 iovss.n653 9.0005
R10022 iovss.n662 iovss.n653 9.0005
R10023 iovss.n719 iovss.n653 9.0005
R10024 iovss.n661 iovss.n653 9.0005
R10025 iovss.n722 iovss.n653 9.0005
R10026 iovss.n660 iovss.n653 9.0005
R10027 iovss.n724 iovss.n653 9.0005
R10028 iovss.n659 iovss.n653 9.0005
R10029 iovss.n727 iovss.n653 9.0005
R10030 iovss.n658 iovss.n653 9.0005
R10031 iovss.n729 iovss.n653 9.0005
R10032 iovss.n657 iovss.n653 9.0005
R10033 iovss.n731 iovss.n653 9.0005
R10034 iovss.n3246 iovss.n653 9.0005
R10035 iovss.n3249 iovss.n653 9.0005
R10036 iovss.n672 iovss.n637 9.0005
R10037 iovss.n676 iovss.n637 9.0005
R10038 iovss.n671 iovss.n637 9.0005
R10039 iovss.n678 iovss.n637 9.0005
R10040 iovss.n670 iovss.n637 9.0005
R10041 iovss.n681 iovss.n637 9.0005
R10042 iovss.n669 iovss.n637 9.0005
R10043 iovss.n683 iovss.n637 9.0005
R10044 iovss.n668 iovss.n637 9.0005
R10045 iovss.n686 iovss.n637 9.0005
R10046 iovss.n667 iovss.n637 9.0005
R10047 iovss.n688 iovss.n637 9.0005
R10048 iovss.n666 iovss.n637 9.0005
R10049 iovss.n691 iovss.n637 9.0005
R10050 iovss.n665 iovss.n637 9.0005
R10051 iovss.n710 iovss.n637 9.0005
R10052 iovss.n664 iovss.n637 9.0005
R10053 iovss.n712 iovss.n637 9.0005
R10054 iovss.n3251 iovss.n637 9.0005
R10055 iovss.n714 iovss.n637 9.0005
R10056 iovss.n663 iovss.n637 9.0005
R10057 iovss.n717 iovss.n637 9.0005
R10058 iovss.n662 iovss.n637 9.0005
R10059 iovss.n719 iovss.n637 9.0005
R10060 iovss.n661 iovss.n637 9.0005
R10061 iovss.n722 iovss.n637 9.0005
R10062 iovss.n660 iovss.n637 9.0005
R10063 iovss.n724 iovss.n637 9.0005
R10064 iovss.n659 iovss.n637 9.0005
R10065 iovss.n727 iovss.n637 9.0005
R10066 iovss.n658 iovss.n637 9.0005
R10067 iovss.n729 iovss.n637 9.0005
R10068 iovss.n657 iovss.n637 9.0005
R10069 iovss.n731 iovss.n637 9.0005
R10070 iovss.n3246 iovss.n637 9.0005
R10071 iovss.n3249 iovss.n637 9.0005
R10072 iovss.n672 iovss.n654 9.0005
R10073 iovss.n676 iovss.n654 9.0005
R10074 iovss.n671 iovss.n654 9.0005
R10075 iovss.n678 iovss.n654 9.0005
R10076 iovss.n670 iovss.n654 9.0005
R10077 iovss.n681 iovss.n654 9.0005
R10078 iovss.n669 iovss.n654 9.0005
R10079 iovss.n683 iovss.n654 9.0005
R10080 iovss.n668 iovss.n654 9.0005
R10081 iovss.n686 iovss.n654 9.0005
R10082 iovss.n667 iovss.n654 9.0005
R10083 iovss.n688 iovss.n654 9.0005
R10084 iovss.n666 iovss.n654 9.0005
R10085 iovss.n691 iovss.n654 9.0005
R10086 iovss.n665 iovss.n654 9.0005
R10087 iovss.n710 iovss.n654 9.0005
R10088 iovss.n664 iovss.n654 9.0005
R10089 iovss.n712 iovss.n654 9.0005
R10090 iovss.n3251 iovss.n654 9.0005
R10091 iovss.n714 iovss.n654 9.0005
R10092 iovss.n663 iovss.n654 9.0005
R10093 iovss.n717 iovss.n654 9.0005
R10094 iovss.n662 iovss.n654 9.0005
R10095 iovss.n719 iovss.n654 9.0005
R10096 iovss.n661 iovss.n654 9.0005
R10097 iovss.n722 iovss.n654 9.0005
R10098 iovss.n660 iovss.n654 9.0005
R10099 iovss.n724 iovss.n654 9.0005
R10100 iovss.n659 iovss.n654 9.0005
R10101 iovss.n727 iovss.n654 9.0005
R10102 iovss.n658 iovss.n654 9.0005
R10103 iovss.n729 iovss.n654 9.0005
R10104 iovss.n657 iovss.n654 9.0005
R10105 iovss.n731 iovss.n654 9.0005
R10106 iovss.n3246 iovss.n654 9.0005
R10107 iovss.n3249 iovss.n654 9.0005
R10108 iovss.n672 iovss.n636 9.0005
R10109 iovss.n676 iovss.n636 9.0005
R10110 iovss.n671 iovss.n636 9.0005
R10111 iovss.n678 iovss.n636 9.0005
R10112 iovss.n670 iovss.n636 9.0005
R10113 iovss.n681 iovss.n636 9.0005
R10114 iovss.n669 iovss.n636 9.0005
R10115 iovss.n683 iovss.n636 9.0005
R10116 iovss.n668 iovss.n636 9.0005
R10117 iovss.n686 iovss.n636 9.0005
R10118 iovss.n667 iovss.n636 9.0005
R10119 iovss.n688 iovss.n636 9.0005
R10120 iovss.n666 iovss.n636 9.0005
R10121 iovss.n691 iovss.n636 9.0005
R10122 iovss.n665 iovss.n636 9.0005
R10123 iovss.n710 iovss.n636 9.0005
R10124 iovss.n664 iovss.n636 9.0005
R10125 iovss.n712 iovss.n636 9.0005
R10126 iovss.n3251 iovss.n636 9.0005
R10127 iovss.n714 iovss.n636 9.0005
R10128 iovss.n663 iovss.n636 9.0005
R10129 iovss.n717 iovss.n636 9.0005
R10130 iovss.n662 iovss.n636 9.0005
R10131 iovss.n719 iovss.n636 9.0005
R10132 iovss.n661 iovss.n636 9.0005
R10133 iovss.n722 iovss.n636 9.0005
R10134 iovss.n660 iovss.n636 9.0005
R10135 iovss.n724 iovss.n636 9.0005
R10136 iovss.n659 iovss.n636 9.0005
R10137 iovss.n727 iovss.n636 9.0005
R10138 iovss.n658 iovss.n636 9.0005
R10139 iovss.n729 iovss.n636 9.0005
R10140 iovss.n657 iovss.n636 9.0005
R10141 iovss.n731 iovss.n636 9.0005
R10142 iovss.n3246 iovss.n636 9.0005
R10143 iovss.n3249 iovss.n636 9.0005
R10144 iovss.n3250 iovss.n672 9.0005
R10145 iovss.n3250 iovss.n676 9.0005
R10146 iovss.n3250 iovss.n671 9.0005
R10147 iovss.n3250 iovss.n678 9.0005
R10148 iovss.n3250 iovss.n670 9.0005
R10149 iovss.n3250 iovss.n681 9.0005
R10150 iovss.n3250 iovss.n669 9.0005
R10151 iovss.n3250 iovss.n683 9.0005
R10152 iovss.n3250 iovss.n668 9.0005
R10153 iovss.n3250 iovss.n686 9.0005
R10154 iovss.n3250 iovss.n667 9.0005
R10155 iovss.n3250 iovss.n688 9.0005
R10156 iovss.n3250 iovss.n666 9.0005
R10157 iovss.n3250 iovss.n691 9.0005
R10158 iovss.n3250 iovss.n665 9.0005
R10159 iovss.n3250 iovss.n710 9.0005
R10160 iovss.n3250 iovss.n664 9.0005
R10161 iovss.n3250 iovss.n712 9.0005
R10162 iovss.n3251 iovss.n3250 9.0005
R10163 iovss.n3250 iovss.n714 9.0005
R10164 iovss.n3250 iovss.n663 9.0005
R10165 iovss.n3250 iovss.n717 9.0005
R10166 iovss.n3250 iovss.n662 9.0005
R10167 iovss.n3250 iovss.n719 9.0005
R10168 iovss.n3250 iovss.n661 9.0005
R10169 iovss.n3250 iovss.n722 9.0005
R10170 iovss.n3250 iovss.n660 9.0005
R10171 iovss.n3250 iovss.n724 9.0005
R10172 iovss.n3250 iovss.n659 9.0005
R10173 iovss.n3250 iovss.n727 9.0005
R10174 iovss.n3250 iovss.n658 9.0005
R10175 iovss.n3250 iovss.n729 9.0005
R10176 iovss.n3250 iovss.n657 9.0005
R10177 iovss.n3250 iovss.n731 9.0005
R10178 iovss.n3250 iovss.n3249 9.0005
R10179 iovss.n3144 iovss.n892 9.0005
R10180 iovss.n3146 iovss.n892 9.0005
R10181 iovss.n3146 iovss.n894 9.0005
R10182 iovss.n3146 iovss.n891 9.0005
R10183 iovss.n3146 iovss.n896 9.0005
R10184 iovss.n3146 iovss.n890 9.0005
R10185 iovss.n3146 iovss.n898 9.0005
R10186 iovss.n3146 iovss.n889 9.0005
R10187 iovss.n3146 iovss.n900 9.0005
R10188 iovss.n3146 iovss.n888 9.0005
R10189 iovss.n3146 iovss.n902 9.0005
R10190 iovss.n3146 iovss.n887 9.0005
R10191 iovss.n3145 iovss.n3144 9.0005
R10192 iovss.n3146 iovss.n3145 9.0005
R10193 iovss.n913 iovss.n907 9.0005
R10194 iovss.n3136 iovss.n913 9.0005
R10195 iovss.n3136 iovss.n915 9.0005
R10196 iovss.n919 iovss.n907 9.0005
R10197 iovss.n3136 iovss.n919 9.0005
R10198 iovss.n3136 iovss.n911 9.0005
R10199 iovss.n1198 iovss.n922 9.0005
R10200 iovss.n3136 iovss.n922 9.0005
R10201 iovss.n910 iovss.n907 9.0005
R10202 iovss.n3136 iovss.n910 9.0005
R10203 iovss.n924 iovss.n907 9.0005
R10204 iovss.n3136 iovss.n924 9.0005
R10205 iovss.n909 iovss.n907 9.0005
R10206 iovss.n3136 iovss.n909 9.0005
R10207 iovss.n3136 iovss.n3135 9.0005
R10208 iovss.n3136 iovss.n908 9.0005
R10209 iovss.n3137 iovss.n907 9.0005
R10210 iovss.n3137 iovss.n3136 9.0005
R10211 iovss.n949 iovss.n938 9.0005
R10212 iovss.n3130 iovss.n938 9.0005
R10213 iovss.n3130 iovss.n940 9.0005
R10214 iovss.n3130 iovss.n937 9.0005
R10215 iovss.n3130 iovss.n942 9.0005
R10216 iovss.n3130 iovss.n936 9.0005
R10217 iovss.n3130 iovss.n944 9.0005
R10218 iovss.n3130 iovss.n935 9.0005
R10219 iovss.n3130 iovss.n3129 9.0005
R10220 iovss.n3130 iovss.n934 9.0005
R10221 iovss.n3131 iovss.n3130 9.0005
R10222 iovss.n3130 iovss.n933 9.0005
R10223 iovss.n949 iovss.n905 9.0005
R10224 iovss.n3130 iovss.n905 9.0005
R10225 iovss.n46 iovss 7.94638
R10226 iovss.t2 iovss.n1350 5.66717
R10227 iovss.n2757 iovss.t2 5.66717
R10228 iovss.t2 iovss.n1379 5.66717
R10229 iovss.t2 iovss.n1376 5.66717
R10230 iovss.t2 iovss.n1384 5.66717
R10231 iovss.t2 iovss.n1374 5.66717
R10232 iovss.t2 iovss.n1386 5.66717
R10233 iovss.t2 iovss.n1373 5.66717
R10234 iovss.t2 iovss.n1388 5.66717
R10235 iovss.t2 iovss.n1371 5.66717
R10236 iovss.t2 iovss.n1390 5.66717
R10237 iovss.t2 iovss.n1369 5.66717
R10238 iovss.t2 iovss.n1391 5.66717
R10239 iovss.t2 iovss.n1367 5.66717
R10240 iovss.t2 iovss.n1393 5.66717
R10241 iovss.t2 iovss.n1365 5.66717
R10242 iovss.t2 iovss.n1394 5.66717
R10243 iovss.t2 iovss.n1363 5.66717
R10244 iovss.t2 iovss.n1396 5.66717
R10245 iovss.t2 iovss.n1361 5.66717
R10246 iovss.t2 iovss.n1398 5.66717
R10247 iovss.t2 iovss.n1360 5.66717
R10248 iovss.t2 iovss.n1400 5.66717
R10249 iovss.t2 iovss.n1358 5.66717
R10250 iovss.t2 iovss.n1402 5.66717
R10251 iovss.t2 iovss.n1356 5.66717
R10252 iovss.t2 iovss.n1403 5.66717
R10253 iovss.t2 iovss.n1354 5.66717
R10254 iovss.t2 iovss.n1405 5.66717
R10255 iovss.t2 iovss.n1352 5.66717
R10256 iovss.t2 iovss.n1407 5.66717
R10257 iovss.t0 iovss.n1278 5.66717
R10258 iovss.t0 iovss.n1276 5.66717
R10259 iovss.t0 iovss.n1279 5.66717
R10260 iovss.t0 iovss.n1274 5.66717
R10261 iovss.t0 iovss.n1281 5.66717
R10262 iovss.t0 iovss.n1272 5.66717
R10263 iovss.t0 iovss.n1283 5.66717
R10264 iovss.t0 iovss.n1271 5.66717
R10265 iovss.t0 iovss.n1286 5.66717
R10266 iovss.t0 iovss.n1269 5.66717
R10267 iovss.t0 iovss.n1288 5.66717
R10268 iovss.t0 iovss.n1267 5.66717
R10269 iovss.t0 iovss.n1289 5.66717
R10270 iovss.t0 iovss.n1265 5.66717
R10271 iovss.t0 iovss.n1291 5.66717
R10272 iovss.t0 iovss.n1263 5.66717
R10273 iovss.t0 iovss.n1292 5.66717
R10274 iovss.t0 iovss.n1261 5.66717
R10275 iovss.t0 iovss.n1294 5.66717
R10276 iovss.t0 iovss.n1259 5.66717
R10277 iovss.t0 iovss.n1296 5.66717
R10278 iovss.t0 iovss.n1258 5.66717
R10279 iovss.t0 iovss.n1298 5.66717
R10280 iovss.t0 iovss.n1256 5.66717
R10281 iovss.t0 iovss.n1300 5.66717
R10282 iovss.t0 iovss.n1254 5.66717
R10283 iovss.t0 iovss.n1301 5.66717
R10284 iovss.t0 iovss.n1252 5.66717
R10285 iovss.t0 iovss.n1303 5.66717
R10286 iovss.t0 iovss.n1250 5.66717
R10287 iovss.t0 iovss.n2894 5.66717
R10288 iovss.n1731 iovss.n303 4.50058
R10289 iovss.n1803 iovss.n303 4.50058
R10290 iovss.n1805 iovss.n303 4.50058
R10291 iovss.n1808 iovss.n303 4.50058
R10292 iovss.n1810 iovss.n303 4.50058
R10293 iovss.n1813 iovss.n303 4.50058
R10294 iovss.n1815 iovss.n303 4.50058
R10295 iovss.n1818 iovss.n303 4.50058
R10296 iovss.n1820 iovss.n303 4.50058
R10297 iovss.n1823 iovss.n303 4.50058
R10298 iovss.n1825 iovss.n303 4.50058
R10299 iovss.n1828 iovss.n303 4.50058
R10300 iovss.n1831 iovss.n303 4.50058
R10301 iovss.n1833 iovss.n303 4.50058
R10302 iovss.n1836 iovss.n303 4.50058
R10303 iovss.n1838 iovss.n303 4.50058
R10304 iovss.n1843 iovss.n303 4.50058
R10305 iovss.n1842 iovss.n303 4.50058
R10306 iovss.n1800 iovss.n1732 4.50058
R10307 iovss.n1806 iovss.n1732 4.50058
R10308 iovss.n1811 iovss.n1732 4.50058
R10309 iovss.n1816 iovss.n1732 4.50058
R10310 iovss.n1821 iovss.n1732 4.50058
R10311 iovss.n1826 iovss.n1732 4.50058
R10312 iovss.n1829 iovss.n1732 4.50058
R10313 iovss.n1834 iovss.n1732 4.50058
R10314 iovss.n1839 iovss.n1732 4.50058
R10315 iovss.n1869 iovss.n1732 4.50058
R10316 iovss.n1917 iovss.n673 4.50058
R10317 iovss.n1959 iovss.n673 4.50058
R10318 iovss.n2096 iovss.n673 4.50058
R10319 iovss.n2099 iovss.n673 4.50058
R10320 iovss.n2102 iovss.n673 4.50058
R10321 iovss.n2105 iovss.n673 4.50058
R10322 iovss.n2107 iovss.n673 4.50058
R10323 iovss.n2110 iovss.n673 4.50058
R10324 iovss.n2112 iovss.n673 4.50058
R10325 iovss.n2115 iovss.n673 4.50058
R10326 iovss.n2117 iovss.n673 4.50058
R10327 iovss.n2122 iovss.n673 4.50058
R10328 iovss.n2127 iovss.n673 4.50058
R10329 iovss.n2158 iovss.n673 4.50058
R10330 iovss.n2094 iovss.n1918 4.50058
R10331 iovss.n2097 iovss.n1918 4.50058
R10332 iovss.n2103 iovss.n1918 4.50058
R10333 iovss.n2108 iovss.n1918 4.50058
R10334 iovss.n2113 iovss.n1918 4.50058
R10335 iovss.n2118 iovss.n1918 4.50058
R10336 iovss.n2120 iovss.n1918 4.50058
R10337 iovss.n2123 iovss.n1918 4.50058
R10338 iovss.n2125 iovss.n1918 4.50058
R10339 iovss.n2128 iovss.n1918 4.50058
R10340 iovss.n2130 iovss.n1918 4.50058
R10341 iovss.n2159 iovss.n1918 4.50058
R10342 iovss.n2242 iovss.n1944 4.50058
R10343 iovss.n3076 iovss.n2901 4.50058
R10344 iovss.n3097 iovss.n3096 4.50058
R10345 iovss.n3094 iovss.n1108 4.50058
R10346 iovss.n1106 iovss.n1105 4.50058
R10347 iovss.n3112 iovss.n961 4.50058
R10348 iovss.n1568 iovss.n220 4.50058
R10349 iovss.n1570 iovss.n220 4.50058
R10350 iovss.n1572 iovss.n220 4.50058
R10351 iovss.n1574 iovss.n220 4.50058
R10352 iovss.n1576 iovss.n220 4.50058
R10353 iovss.n1578 iovss.n220 4.50058
R10354 iovss.n1580 iovss.n220 4.50058
R10355 iovss.n1582 iovss.n220 4.50058
R10356 iovss.n1584 iovss.n220 4.50058
R10357 iovss.n1586 iovss.n220 4.50058
R10358 iovss.n1588 iovss.n220 4.50058
R10359 iovss.n1590 iovss.n220 4.50058
R10360 iovss.n1592 iovss.n220 4.50058
R10361 iovss.n1594 iovss.n220 4.50058
R10362 iovss.n1597 iovss.n220 4.50058
R10363 iovss.n1625 iovss.n220 4.50058
R10364 iovss.n2393 iovss.n2392 4.50058
R10365 iovss.n2393 iovss.n2391 4.50058
R10366 iovss.n2393 iovss.n2390 4.50058
R10367 iovss.n2393 iovss.n2389 4.50058
R10368 iovss.n2393 iovss.n2388 4.50058
R10369 iovss.n2393 iovss.n2387 4.50058
R10370 iovss.n2393 iovss.n2386 4.50058
R10371 iovss.n2393 iovss.n2385 4.50058
R10372 iovss.n2393 iovss.n2384 4.50058
R10373 iovss.n2393 iovss.n2383 4.50058
R10374 iovss.n2393 iovss.n2382 4.50058
R10375 iovss.n2393 iovss.n1626 4.50058
R10376 iovss.n2397 iovss.n1550 4.50058
R10377 iovss.n2897 iovss.n1224 4.50058
R10378 iovss.n2752 iovss.n2711 4.50058
R10379 iovss.n2718 iovss.n2716 4.50058
R10380 iovss.n2776 iovss.n1310 4.50058
R10381 iovss.n221 iovss.n172 4.50058
R10382 iovss.n223 iovss.n172 4.50058
R10383 iovss.n225 iovss.n172 4.50058
R10384 iovss.n227 iovss.n172 4.50058
R10385 iovss.n229 iovss.n172 4.50058
R10386 iovss.n231 iovss.n172 4.50058
R10387 iovss.n233 iovss.n172 4.50058
R10388 iovss.n235 iovss.n172 4.50058
R10389 iovss.n185 iovss.n172 4.50058
R10390 iovss.n238 iovss.n172 4.50058
R10391 iovss.n240 iovss.n172 4.50058
R10392 iovss.n242 iovss.n172 4.50058
R10393 iovss.n244 iovss.n172 4.50058
R10394 iovss.n246 iovss.n172 4.50058
R10395 iovss.n249 iovss.n172 4.50058
R10396 iovss.n252 iovss.n172 4.50058
R10397 iovss.n3426 iovss.n3425 4.50058
R10398 iovss.n3426 iovss.n3424 4.50058
R10399 iovss.n3426 iovss.n3423 4.50058
R10400 iovss.n3426 iovss.n3422 4.50058
R10401 iovss.n3426 iovss.n175 4.50058
R10402 iovss.n3426 iovss.n3421 4.50058
R10403 iovss.n3426 iovss.n3420 4.50058
R10404 iovss.n3426 iovss.n3419 4.50058
R10405 iovss.n3426 iovss.n3418 4.50058
R10406 iovss.n3426 iovss.n3417 4.50058
R10407 iovss.n3426 iovss.n3416 4.50058
R10408 iovss.n304 iovss.n275 4.50058
R10409 iovss.n307 iovss.n275 4.50058
R10410 iovss.n310 iovss.n275 4.50058
R10411 iovss.n313 iovss.n275 4.50058
R10412 iovss.n316 iovss.n275 4.50058
R10413 iovss.n319 iovss.n275 4.50058
R10414 iovss.n321 iovss.n275 4.50058
R10415 iovss.n323 iovss.n275 4.50058
R10416 iovss.n325 iovss.n275 4.50058
R10417 iovss.n327 iovss.n275 4.50058
R10418 iovss.n329 iovss.n275 4.50058
R10419 iovss.n3386 iovss.n275 4.50058
R10420 iovss.n3391 iovss.n265 4.50058
R10421 iovss.n3391 iovss.n349 4.50058
R10422 iovss.n3391 iovss.n348 4.50058
R10423 iovss.n3391 iovss.n347 4.50058
R10424 iovss.n3391 iovss.n346 4.50058
R10425 iovss.n3391 iovss.n345 4.50058
R10426 iovss.n3391 iovss.n344 4.50058
R10427 iovss.n3391 iovss.n343 4.50058
R10428 iovss.n3391 iovss.n342 4.50058
R10429 iovss.n3391 iovss.n341 4.50058
R10430 iovss.n3391 iovss.n340 4.50058
R10431 iovss.n3391 iovss.n339 4.50058
R10432 iovss.n3391 iovss.n338 4.50058
R10433 iovss.n3391 iovss.n337 4.50058
R10434 iovss.n3393 iovss.n286 4.50058
R10435 iovss.n674 iovss.n632 4.50058
R10436 iovss.n677 iovss.n632 4.50058
R10437 iovss.n679 iovss.n632 4.50058
R10438 iovss.n682 iovss.n632 4.50058
R10439 iovss.n684 iovss.n632 4.50058
R10440 iovss.n687 iovss.n632 4.50058
R10441 iovss.n689 iovss.n632 4.50058
R10442 iovss.n692 iovss.n632 4.50058
R10443 iovss.n645 iovss.n632 4.50058
R10444 iovss.n713 iovss.n632 4.50058
R10445 iovss.n715 iovss.n632 4.50058
R10446 iovss.n720 iovss.n632 4.50058
R10447 iovss.n725 iovss.n632 4.50058
R10448 iovss.n766 iovss.n632 4.50058
R10449 iovss.n675 iovss.n646 4.50058
R10450 iovss.n680 iovss.n646 4.50058
R10451 iovss.n685 iovss.n646 4.50058
R10452 iovss.n690 iovss.n646 4.50058
R10453 iovss.n711 iovss.n646 4.50058
R10454 iovss.n716 iovss.n646 4.50058
R10455 iovss.n718 iovss.n646 4.50058
R10456 iovss.n721 iovss.n646 4.50058
R10457 iovss.n723 iovss.n646 4.50058
R10458 iovss.n726 iovss.n646 4.50058
R10459 iovss.n728 iovss.n646 4.50058
R10460 iovss.n730 iovss.n646 4.50058
R10461 iovss.n3250 iovss.n656 4.50058
R10462 iovss.n917 iovss.n912 4.50058
R10463 iovss.n2076 iovss.n2034 4.5005
R10464 iovss.n2075 iovss.n2073 4.5005
R10465 iovss.n2037 iovss.n2036 4.5005
R10466 iovss.n2069 iovss.n2068 4.5005
R10467 iovss.n2066 iovss.n2042 4.5005
R10468 iovss.n2064 iovss.n2062 4.5005
R10469 iovss.n2045 iovss.n2044 4.5005
R10470 iovss.n2058 iovss.n2057 4.5005
R10471 iovss.n2055 iovss.n2053 4.5005
R10472 iovss.n1506 iovss.n1503 4.5005
R10473 iovss.n2539 iovss.n2538 4.5005
R10474 iovss.n1507 iovss.n1505 4.5005
R10475 iovss.n2534 iovss.n2533 4.5005
R10476 iovss.n2531 iovss.n1513 4.5005
R10477 iovss.n2529 iovss.n2527 4.5005
R10478 iovss.n1516 iovss.n1515 4.5005
R10479 iovss.n2523 iovss.n2522 4.5005
R10480 iovss.n2520 iovss.n1522 4.5005
R10481 iovss.n2519 iovss.n2517 4.5005
R10482 iovss.n1524 iovss.n1523 4.5005
R10483 iovss.n2513 iovss.n2512 4.5005
R10484 iovss.n1531 iovss.n1530 4.5005
R10485 iovss.n2492 iovss.n2491 4.5005
R10486 iovss.n2405 iovss.n2404 4.5005
R10487 iovss.n2487 iovss.n2486 4.5005
R10488 iovss.n2412 iovss.n2411 4.5005
R10489 iovss.n2468 iovss.n2467 4.5005
R10490 iovss.n2429 iovss.n2428 4.5005
R10491 iovss.n2463 iovss.n2462 4.5005
R10492 iovss.n2437 iovss.n2436 4.5005
R10493 iovss.n1433 iovss.n1432 4.5005
R10494 iovss.n2589 iovss.n2588 4.5005
R10495 iovss.n1427 iovss.n1414 4.5005
R10496 iovss.n2596 iovss.n2595 4.5005
R10497 iovss.n1428 iovss.n1426 4.5005
R10498 iovss.n1426 iovss.n1425 4.5005
R10499 iovss.n2597 iovss.n2596 4.5005
R10500 iovss.n2580 iovss.n1414 4.5005
R10501 iovss.n2588 iovss.n2587 4.5005
R10502 iovss.n1437 iovss.n1433 4.5005
R10503 iovss.n2453 iovss.n2437 4.5005
R10504 iovss.n2462 iovss.n2461 4.5005
R10505 iovss.n2444 iovss.n2428 4.5005
R10506 iovss.n2469 iovss.n2468 4.5005
R10507 iovss.n2477 iovss.n2412 4.5005
R10508 iovss.n2486 iovss.n2485 4.5005
R10509 iovss.n2419 iovss.n2404 4.5005
R10510 iovss.n2493 iovss.n2492 4.5005
R10511 iovss.n2501 iovss.n1531 4.5005
R10512 iovss.n2512 iovss.n2511 4.5005
R10513 iovss.n1537 iovss.n1523 4.5005
R10514 iovss.n2519 iovss.n2518 4.5005
R10515 iovss.n2520 iovss.n1463 4.5005
R10516 iovss.n2522 iovss.n2521 4.5005
R10517 iovss.n1515 iovss.n1514 4.5005
R10518 iovss.n2529 iovss.n2528 4.5005
R10519 iovss.n2531 iovss.n2530 4.5005
R10520 iovss.n2533 iovss.n2532 4.5005
R10521 iovss.n1505 iovss.n1504 4.5005
R10522 iovss.n2540 iovss.n2539 4.5005
R10523 iovss.n1985 iovss.n1503 4.5005
R10524 iovss.n2055 iovss.n2054 4.5005
R10525 iovss.n2057 iovss.n2056 4.5005
R10526 iovss.n2044 iovss.n2043 4.5005
R10527 iovss.n2064 iovss.n2063 4.5005
R10528 iovss.n2066 iovss.n2065 4.5005
R10529 iovss.n2068 iovss.n2067 4.5005
R10530 iovss.n2036 iovss.n2035 4.5005
R10531 iovss.n2075 iovss.n2074 4.5005
R10532 iovss.n2077 iovss.n2076 4.5005
R10533 iovss.n171 iovss.n169 4.50042
R10534 iovss.n171 iovss.n168 4.50042
R10535 iovss.n171 iovss.n167 4.50042
R10536 iovss.n171 iovss.n166 4.50042
R10537 iovss.n171 iovss.n165 4.50042
R10538 iovss.n171 iovss.n164 4.50042
R10539 iovss.n171 iovss.n119 4.50042
R10540 iovss.n2356 iovss.n2355 4.50042
R10541 iovss.n2355 iovss.n1676 4.50042
R10542 iovss.n2355 iovss.n1675 4.50042
R10543 iovss.n2355 iovss.n1674 4.50042
R10544 iovss.n2355 iovss.n1673 4.50042
R10545 iovss.n2355 iovss.n1672 4.50042
R10546 iovss.n2355 iovss.n1671 4.50042
R10547 iovss.n2355 iovss.n1670 4.50042
R10548 iovss.n2355 iovss.n1669 4.50042
R10549 iovss.n2355 iovss.n1668 4.50042
R10550 iovss.n2355 iovss.n1667 4.50042
R10551 iovss.n2355 iovss.n1666 4.50042
R10552 iovss.n2355 iovss.n1665 4.50042
R10553 iovss.n2355 iovss.n1664 4.50042
R10554 iovss.n2355 iovss.n1663 4.50042
R10555 iovss.n2355 iovss.n1662 4.50042
R10556 iovss.n2355 iovss.n1661 4.50042
R10557 iovss.n2355 iovss.n1660 4.50042
R10558 iovss.n2355 iovss.n1659 4.50042
R10559 iovss.n2355 iovss.n1658 4.50042
R10560 iovss.n2355 iovss.n1657 4.50042
R10561 iovss.n2355 iovss.n1656 4.50042
R10562 iovss.n2355 iovss.n1655 4.50042
R10563 iovss.n2355 iovss.n1654 4.50042
R10564 iovss.n2355 iovss.n1650 4.50042
R10565 iovss.n2355 iovss.n1549 4.50042
R10566 iovss.n2024 iovss.n1973 4.50042
R10567 iovss.n2079 iovss.n1999 4.50042
R10568 iovss.n1999 iovss.n1998 4.50042
R10569 iovss.n2080 iovss.n1997 4.50042
R10570 iovss.n2558 iovss.n2557 4.50042
R10571 iovss.n2555 iovss.n2553 4.50042
R10572 iovss.n2558 iovss.n1449 4.50042
R10573 iovss.n2556 iovss.n2555 4.50042
R10574 iovss.n2290 iovss.n2289 4.50042
R10575 iovss.n1783 iovss.n1782 4.50042
R10576 iovss.n1868 iovss.n1844 4.50042
R10577 iovss.n1783 iovss.n1781 4.50042
R10578 iovss.n1868 iovss.n1845 4.50042
R10579 iovss.n1783 iovss.n1780 4.50042
R10580 iovss.n1868 iovss.n1846 4.50042
R10581 iovss.n1783 iovss.n1779 4.50042
R10582 iovss.n1868 iovss.n1847 4.50042
R10583 iovss.n1783 iovss.n1778 4.50042
R10584 iovss.n1868 iovss.n1848 4.50042
R10585 iovss.n1783 iovss.n1777 4.50042
R10586 iovss.n1868 iovss.n1849 4.50042
R10587 iovss.n1783 iovss.n1776 4.50042
R10588 iovss.n1868 iovss.n1850 4.50042
R10589 iovss.n1783 iovss.n1775 4.50042
R10590 iovss.n1868 iovss.n1851 4.50042
R10591 iovss.n1783 iovss.n1774 4.50042
R10592 iovss.n1868 iovss.n1852 4.50042
R10593 iovss.n1783 iovss.n1773 4.50042
R10594 iovss.n1868 iovss.n1853 4.50042
R10595 iovss.n1783 iovss.n1772 4.50042
R10596 iovss.n1868 iovss.n1854 4.50042
R10597 iovss.n1783 iovss.n1771 4.50042
R10598 iovss.n1868 iovss.n1855 4.50042
R10599 iovss.n1783 iovss.n1770 4.50042
R10600 iovss.n1868 iovss.n1856 4.50042
R10601 iovss.n1783 iovss.n1769 4.50042
R10602 iovss.n1868 iovss.n1857 4.50042
R10603 iovss.n1783 iovss.n1768 4.50042
R10604 iovss.n1868 iovss.n1858 4.50042
R10605 iovss.n1783 iovss.n1767 4.50042
R10606 iovss.n1868 iovss.n1859 4.50042
R10607 iovss.n1783 iovss.n1766 4.50042
R10608 iovss.n1868 iovss.n1860 4.50042
R10609 iovss.n1783 iovss.n1765 4.50042
R10610 iovss.n1868 iovss.n1861 4.50042
R10611 iovss.n1783 iovss.n1764 4.50042
R10612 iovss.n1868 iovss.n1862 4.50042
R10613 iovss.n1783 iovss.n1763 4.50042
R10614 iovss.n1868 iovss.n1863 4.50042
R10615 iovss.n1783 iovss.n1762 4.50042
R10616 iovss.n1868 iovss.n1864 4.50042
R10617 iovss.n1783 iovss.n1761 4.50042
R10618 iovss.n1868 iovss.n1865 4.50042
R10619 iovss.n1783 iovss.n1760 4.50042
R10620 iovss.n1868 iovss.n1866 4.50042
R10621 iovss.n1783 iovss.n1759 4.50042
R10622 iovss.n1868 iovss.n1867 4.50042
R10623 iovss.n1783 iovss.n1758 4.50042
R10624 iovss.n1868 iovss.n1757 4.50042
R10625 iovss.n2240 iovss.n2215 4.50042
R10626 iovss.n2157 iovss.n2156 4.50042
R10627 iovss.n2240 iovss.n2216 4.50042
R10628 iovss.n2157 iovss.n2155 4.50042
R10629 iovss.n2240 iovss.n2217 4.50042
R10630 iovss.n2157 iovss.n2154 4.50042
R10631 iovss.n2240 iovss.n2218 4.50042
R10632 iovss.n2157 iovss.n2153 4.50042
R10633 iovss.n2240 iovss.n2219 4.50042
R10634 iovss.n2157 iovss.n2152 4.50042
R10635 iovss.n2240 iovss.n2220 4.50042
R10636 iovss.n2157 iovss.n2151 4.50042
R10637 iovss.n2240 iovss.n2221 4.50042
R10638 iovss.n2157 iovss.n2150 4.50042
R10639 iovss.n2240 iovss.n2222 4.50042
R10640 iovss.n2157 iovss.n2149 4.50042
R10641 iovss.n2240 iovss.n2223 4.50042
R10642 iovss.n2157 iovss.n2148 4.50042
R10643 iovss.n2240 iovss.n2224 4.50042
R10644 iovss.n2157 iovss.n2147 4.50042
R10645 iovss.n2240 iovss.n2225 4.50042
R10646 iovss.n2157 iovss.n2146 4.50042
R10647 iovss.n2240 iovss.n2226 4.50042
R10648 iovss.n2157 iovss.n2145 4.50042
R10649 iovss.n2240 iovss.n2227 4.50042
R10650 iovss.n2157 iovss.n2144 4.50042
R10651 iovss.n2240 iovss.n2228 4.50042
R10652 iovss.n2157 iovss.n2143 4.50042
R10653 iovss.n2240 iovss.n2229 4.50042
R10654 iovss.n2157 iovss.n2142 4.50042
R10655 iovss.n2240 iovss.n2230 4.50042
R10656 iovss.n2157 iovss.n2141 4.50042
R10657 iovss.n2240 iovss.n2231 4.50042
R10658 iovss.n2157 iovss.n2140 4.50042
R10659 iovss.n2240 iovss.n2232 4.50042
R10660 iovss.n2157 iovss.n2139 4.50042
R10661 iovss.n2240 iovss.n2233 4.50042
R10662 iovss.n2157 iovss.n2138 4.50042
R10663 iovss.n2240 iovss.n2234 4.50042
R10664 iovss.n2157 iovss.n2137 4.50042
R10665 iovss.n2240 iovss.n2235 4.50042
R10666 iovss.n2157 iovss.n2136 4.50042
R10667 iovss.n2240 iovss.n2236 4.50042
R10668 iovss.n2157 iovss.n2135 4.50042
R10669 iovss.n2240 iovss.n2237 4.50042
R10670 iovss.n2157 iovss.n2134 4.50042
R10671 iovss.n2240 iovss.n2238 4.50042
R10672 iovss.n2157 iovss.n2133 4.50042
R10673 iovss.n2240 iovss.n2239 4.50042
R10674 iovss.n2157 iovss.n2132 4.50042
R10675 iovss.n2240 iovss.n1943 4.50042
R10676 iovss.n615 iovss.n614 4.50042
R10677 iovss.n518 iovss.n511 4.50042
R10678 iovss.n499 iovss.n489 4.50042
R10679 iovss.n518 iovss.n512 4.50042
R10680 iovss.n501 iovss.n489 4.50042
R10681 iovss.n518 iovss.n513 4.50042
R10682 iovss.n503 iovss.n489 4.50042
R10683 iovss.n518 iovss.n514 4.50042
R10684 iovss.n505 iovss.n489 4.50042
R10685 iovss.n518 iovss.n515 4.50042
R10686 iovss.n507 iovss.n489 4.50042
R10687 iovss.n518 iovss.n516 4.50042
R10688 iovss.n509 iovss.n489 4.50042
R10689 iovss.n518 iovss.n517 4.50042
R10690 iovss.n520 iovss.n489 4.50042
R10691 iovss.n3333 iovss.n360 4.50042
R10692 iovss.n409 iovss.n402 4.50042
R10693 iovss.n390 iovss.n362 4.50042
R10694 iovss.n409 iovss.n403 4.50042
R10695 iovss.n392 iovss.n362 4.50042
R10696 iovss.n409 iovss.n404 4.50042
R10697 iovss.n394 iovss.n362 4.50042
R10698 iovss.n409 iovss.n405 4.50042
R10699 iovss.n396 iovss.n362 4.50042
R10700 iovss.n409 iovss.n406 4.50042
R10701 iovss.n398 iovss.n362 4.50042
R10702 iovss.n409 iovss.n407 4.50042
R10703 iovss.n400 iovss.n362 4.50042
R10704 iovss.n409 iovss.n408 4.50042
R10705 iovss.n411 iovss.n362 4.50042
R10706 iovss.n149 iovss.n101 4.50042
R10707 iovss.n103 iovss.n102 4.50042
R10708 iovss.n101 iovss.n95 4.50042
R10709 iovss.n101 iovss.n96 4.50042
R10710 iovss.n101 iovss.n97 4.50042
R10711 iovss.n101 iovss.n98 4.50042
R10712 iovss.n101 iovss.n99 4.50042
R10713 iovss.n101 iovss.n100 4.50042
R10714 iovss.n2381 iovss.n2380 4.50042
R10715 iovss.n2380 iovss.n2379 4.50042
R10716 iovss.n2380 iovss.n2378 4.50042
R10717 iovss.n2380 iovss.n2377 4.50042
R10718 iovss.n2380 iovss.n2376 4.50042
R10719 iovss.n2380 iovss.n2375 4.50042
R10720 iovss.n2380 iovss.n2374 4.50042
R10721 iovss.n2380 iovss.n2373 4.50042
R10722 iovss.n2380 iovss.n2372 4.50042
R10723 iovss.n2380 iovss.n2371 4.50042
R10724 iovss.n2380 iovss.n2370 4.50042
R10725 iovss.n2380 iovss.n2369 4.50042
R10726 iovss.n2380 iovss.n2368 4.50042
R10727 iovss.n2380 iovss.n2367 4.50042
R10728 iovss.n2380 iovss.n2366 4.50042
R10729 iovss.n2380 iovss.n2365 4.50042
R10730 iovss.n2380 iovss.n2364 4.50042
R10731 iovss.n2380 iovss.n2363 4.50042
R10732 iovss.n2380 iovss.n2362 4.50042
R10733 iovss.n2380 iovss.n2361 4.50042
R10734 iovss.n2380 iovss.n2360 4.50042
R10735 iovss.n2380 iovss.n2359 4.50042
R10736 iovss.n2380 iovss.n2358 4.50042
R10737 iovss.n2380 iovss.n2357 4.50042
R10738 iovss.n2380 iovss.n1651 4.50042
R10739 iovss.n2508 iovss.n2507 4.50042
R10740 iovss.n2503 iovss.n2402 4.50042
R10741 iovss.n2508 iovss.n2401 4.50042
R10742 iovss.n2503 iovss.n2502 4.50042
R10743 iovss.n3414 iovss.n263 4.50042
R10744 iovss.n3415 iovss.n203 4.50042
R10745 iovss.n263 iovss.n255 4.50042
R10746 iovss.n203 iovss.n202 4.50042
R10747 iovss.n263 iovss.n256 4.50042
R10748 iovss.n203 iovss.n201 4.50042
R10749 iovss.n263 iovss.n257 4.50042
R10750 iovss.n203 iovss.n200 4.50042
R10751 iovss.n263 iovss.n258 4.50042
R10752 iovss.n203 iovss.n199 4.50042
R10753 iovss.n263 iovss.n259 4.50042
R10754 iovss.n203 iovss.n198 4.50042
R10755 iovss.n263 iovss.n260 4.50042
R10756 iovss.n203 iovss.n197 4.50042
R10757 iovss.n263 iovss.n261 4.50042
R10758 iovss.n203 iovss.n196 4.50042
R10759 iovss.n263 iovss.n262 4.50042
R10760 iovss.n203 iovss.n195 4.50042
R10761 iovss.n263 iovss.n194 4.50042
R10762 iovss.n358 iovss.n335 4.50042
R10763 iovss.n3387 iovss.n336 4.50042
R10764 iovss.n358 iovss.n350 4.50042
R10765 iovss.n3387 iovss.n3385 4.50042
R10766 iovss.n358 iovss.n351 4.50042
R10767 iovss.n3387 iovss.n3384 4.50042
R10768 iovss.n358 iovss.n352 4.50042
R10769 iovss.n3387 iovss.n3383 4.50042
R10770 iovss.n358 iovss.n353 4.50042
R10771 iovss.n3387 iovss.n3382 4.50042
R10772 iovss.n358 iovss.n354 4.50042
R10773 iovss.n3387 iovss.n3381 4.50042
R10774 iovss.n358 iovss.n355 4.50042
R10775 iovss.n3387 iovss.n3380 4.50042
R10776 iovss.n358 iovss.n356 4.50042
R10777 iovss.n3387 iovss.n3379 4.50042
R10778 iovss.n358 iovss.n357 4.50042
R10779 iovss.n3387 iovss.n3378 4.50042
R10780 iovss.n358 iovss.n285 4.50042
R10781 iovss.n742 iovss.n733 4.50042
R10782 iovss.n767 iovss.n765 4.50042
R10783 iovss.n742 iovss.n734 4.50042
R10784 iovss.n767 iovss.n764 4.50042
R10785 iovss.n742 iovss.n735 4.50042
R10786 iovss.n767 iovss.n763 4.50042
R10787 iovss.n742 iovss.n736 4.50042
R10788 iovss.n767 iovss.n762 4.50042
R10789 iovss.n742 iovss.n737 4.50042
R10790 iovss.n767 iovss.n761 4.50042
R10791 iovss.n742 iovss.n738 4.50042
R10792 iovss.n767 iovss.n760 4.50042
R10793 iovss.n742 iovss.n739 4.50042
R10794 iovss.n767 iovss.n759 4.50042
R10795 iovss.n742 iovss.n740 4.50042
R10796 iovss.n767 iovss.n758 4.50042
R10797 iovss.n742 iovss.n741 4.50042
R10798 iovss.n767 iovss.n757 4.50042
R10799 iovss.n742 iovss.n655 4.50042
R10800 iovss.n3254 iovss.n631 4.49965
R10801 iovss.n3254 iovss.n630 4.49965
R10802 iovss.n3254 iovss.n629 4.49965
R10803 iovss.n3254 iovss.n628 4.49965
R10804 iovss.n3254 iovss.n627 4.49965
R10805 iovss.n3254 iovss.n626 4.49965
R10806 iovss.n3254 iovss.n625 4.49965
R10807 iovss.n3254 iovss.n624 4.49965
R10808 iovss.n3254 iovss.n623 4.49965
R10809 iovss.n3254 iovss.n622 4.49965
R10810 iovss.n3254 iovss.n621 4.49965
R10811 iovss.n3254 iovss.n620 4.49965
R10812 iovss.n3254 iovss.n619 4.49965
R10813 iovss.n3254 iovss.n618 4.49965
R10814 iovss.n3254 iovss.n617 4.49965
R10815 iovss.n3254 iovss.n616 4.49965
R10816 iovss.n3255 iovss.n3254 4.49965
R10817 iovss.n3254 iovss.n497 4.49965
R10818 iovss.n539 iovss.n498 4.49965
R10819 iovss.n542 iovss.n498 4.49965
R10820 iovss.n545 iovss.n498 4.49965
R10821 iovss.n548 iovss.n498 4.49965
R10822 iovss.n550 iovss.n498 4.49965
R10823 iovss.n553 iovss.n498 4.49965
R10824 iovss.n556 iovss.n498 4.49965
R10825 iovss.n610 iovss.n498 4.49965
R10826 iovss.n3256 iovss.n498 4.49965
R10827 iovss.n3258 iovss.n519 4.49965
R10828 iovss.n3344 iovss.n379 4.49965
R10829 iovss.n3344 iovss.n378 4.49965
R10830 iovss.n3344 iovss.n377 4.49965
R10831 iovss.n3344 iovss.n376 4.49965
R10832 iovss.n3344 iovss.n375 4.49965
R10833 iovss.n3344 iovss.n374 4.49965
R10834 iovss.n3344 iovss.n372 4.49965
R10835 iovss.n3344 iovss.n371 4.49965
R10836 iovss.n3344 iovss.n370 4.49965
R10837 iovss.n3344 iovss.n369 4.49965
R10838 iovss.n3344 iovss.n368 4.49965
R10839 iovss.n3344 iovss.n367 4.49965
R10840 iovss.n3344 iovss.n366 4.49965
R10841 iovss.n3344 iovss.n365 4.49965
R10842 iovss.n3344 iovss.n364 4.49965
R10843 iovss.n3344 iovss.n363 4.49965
R10844 iovss.n3344 iovss.n361 4.49965
R10845 iovss.n430 iovss.n389 4.49965
R10846 iovss.n433 iovss.n389 4.49965
R10847 iovss.n436 iovss.n389 4.49965
R10848 iovss.n421 iovss.n389 4.49965
R10849 iovss.n438 iovss.n389 4.49965
R10850 iovss.n441 iovss.n389 4.49965
R10851 iovss.n444 iovss.n389 4.49965
R10852 iovss.n447 iovss.n389 4.49965
R10853 iovss.n450 iovss.n389 4.49965
R10854 iovss.n3340 iovss.n389 4.49965
R10855 iovss.n3342 iovss.n410 4.49965
R10856 iovss.n3477 iovss.n3476 4.49965
R10857 iovss.n3476 iovss.n3475 4.49965
R10858 iovss.n3476 iovss.n3474 4.49965
R10859 iovss.n3476 iovss.n3473 4.49965
R10860 iovss.n3476 iovss.n3472 4.49965
R10861 iovss.n3476 iovss.n0 4.49965
R10862 iovss.n50 iovss.n8 4.49965
R10863 iovss.n53 iovss.n8 4.49965
R10864 iovss.n56 iovss.n8 4.49965
R10865 iovss.n3432 iovss.n163 4.49965
R10866 iovss.n3432 iovss.n162 4.49965
R10867 iovss.n3432 iovss.n161 4.49965
R10868 iovss.n3432 iovss.n160 4.49965
R10869 iovss.n3432 iovss.n159 4.49965
R10870 iovss.n3432 iovss.n158 4.49965
R10871 iovss.n3432 iovss.n157 4.49965
R10872 iovss.n3432 iovss.n156 4.49965
R10873 iovss.n3432 iovss.n155 4.49965
R10874 iovss.n3432 iovss.n154 4.49965
R10875 iovss.n3432 iovss.n153 4.49965
R10876 iovss.n3432 iovss.n152 4.49965
R10877 iovss.n3432 iovss.n151 4.49965
R10878 iovss.n3432 iovss.n150 4.49965
R10879 iovss.n3432 iovss.n86 4.49965
R10880 iovss.n170 iovss.n87 4.49965
R10881 iovss.n121 iovss.n87 4.49965
R10882 iovss.n123 iovss.n87 4.49965
R10883 iovss.n125 iovss.n87 4.49965
R10884 iovss.n127 iovss.n87 4.49965
R10885 iovss.n129 iovss.n87 4.49965
R10886 iovss.n131 iovss.n87 4.49965
R10887 iovss.n133 iovss.n87 4.49965
R10888 iovss.n136 iovss.n87 4.49965
R10889 iovss.n139 iovss.n87 4.49965
R10890 iovss.n142 iovss.n87 4.49965
R10891 iovss.n146 iovss.n87 4.49965
R10892 iovss.n148 iovss.n85 4.49965
R10893 iovss.n3433 iovss.n88 4.49965
R10894 iovss.n3105 iovss.n1034 4.49912
R10895 iovss.n3471 iovss.n31 4.4991
R10896 iovss.n31 iovss.n30 4.4991
R10897 iovss.n31 iovss.n29 4.4991
R10898 iovss.n31 iovss.n28 4.4991
R10899 iovss.n35 iovss.n34 4.4991
R10900 iovss.n31 iovss.n27 4.4991
R10901 iovss.n31 iovss.n26 4.4991
R10902 iovss.n44 iovss.n43 4.4991
R10903 iovss.n35 iovss.n33 4.4991
R10904 iovss.n44 iovss.n42 4.4991
R10905 iovss.n44 iovss.n41 4.4991
R10906 iovss.n35 iovss.n32 4.4991
R10907 iovss.n44 iovss.n40 4.4991
R10908 iovss.n44 iovss.n39 4.4991
R10909 iovss.n44 iovss.n15 4.4991
R10910 iovss.n2093 iovss.n1980 4.49741
R10911 iovss.n2093 iovss.n1979 4.49741
R10912 iovss.n2093 iovss.n1978 4.49741
R10913 iovss.n2093 iovss.n1977 4.49741
R10914 iovss.n2093 iovss.n1976 4.49741
R10915 iovss.n2093 iovss.n1975 4.49741
R10916 iovss.n2093 iovss.n1974 4.49741
R10917 iovss.n2093 iovss.n1972 4.49741
R10918 iovss.n2093 iovss.n1971 4.49741
R10919 iovss.n2093 iovss.n1970 4.49741
R10920 iovss.n2093 iovss.n1969 4.49741
R10921 iovss.n2093 iovss.n1968 4.49741
R10922 iovss.n2093 iovss.n1967 4.49741
R10923 iovss.n2093 iovss.n1966 4.49741
R10924 iovss.n2093 iovss.n1965 4.49741
R10925 iovss.n2093 iovss.n1964 4.49741
R10926 iovss.n2093 iovss.n1963 4.49741
R10927 iovss.n2093 iovss.n1962 4.49741
R10928 iovss.n2089 iovss.n1981 4.49741
R10929 iovss.n2089 iovss.n2088 4.49741
R10930 iovss.n2089 iovss.n2087 4.49741
R10931 iovss.n2089 iovss.n2086 4.49741
R10932 iovss.n2089 iovss.n2085 4.49741
R10933 iovss.n2089 iovss.n2084 4.49741
R10934 iovss.n2089 iovss.n2083 4.49741
R10935 iovss.n2089 iovss.n2082 4.49741
R10936 iovss.n2089 iovss.n2081 4.49741
R10937 iovss.n2023 iovss.n1440 4.49741
R10938 iovss.n1541 iovss.n1442 4.49741
R10939 iovss.n1540 iovss.n1445 4.49741
R10940 iovss.n1544 iovss.n1532 4.49741
R10941 iovss.n1993 iovss.n1984 4.49741
R10942 iovss.n1992 iovss.n1446 4.49741
R10943 iovss.n1502 iovss.n1501 4.49741
R10944 iovss.n1502 iovss.n1500 4.49741
R10945 iovss.n1502 iovss.n1499 4.49741
R10946 iovss.n1502 iovss.n1498 4.49741
R10947 iovss.n1502 iovss.n1497 4.49741
R10948 iovss.n1502 iovss.n1496 4.49741
R10949 iovss.n1502 iovss.n1495 4.49741
R10950 iovss.n1502 iovss.n1494 4.49741
R10951 iovss.n1502 iovss.n1493 4.49741
R10952 iovss.n1502 iovss.n1492 4.49741
R10953 iovss.n1502 iovss.n1491 4.49741
R10954 iovss.n1502 iovss.n1490 4.49741
R10955 iovss.n1502 iovss.n1489 4.49741
R10956 iovss.n1502 iovss.n1488 4.49741
R10957 iovss.n1502 iovss.n1487 4.49741
R10958 iovss.n2554 iovss.n1502 4.49741
R10959 iovss.n2552 iovss.n2551 4.49741
R10960 iovss.n2552 iovss.n2550 4.49741
R10961 iovss.n2552 iovss.n2549 4.49741
R10962 iovss.n2552 iovss.n2548 4.49741
R10963 iovss.n2552 iovss.n2547 4.49741
R10964 iovss.n2552 iovss.n2546 4.49741
R10965 iovss.n2552 iovss.n2545 4.49741
R10966 iovss.n2552 iovss.n2544 4.49741
R10967 iovss.n2552 iovss.n2543 4.49741
R10968 iovss.n2552 iovss.n2542 4.49741
R10969 iovss.n2552 iovss.n2541 4.49741
R10970 iovss.n2559 iovss.n1448 4.49741
R10971 iovss.n2563 iovss.n1450 4.49741
R10972 iovss.n2457 iovss.n2398 4.49741
R10973 iovss.n2448 iovss.n2398 4.49741
R10974 iovss.n2440 iovss.n2398 4.49741
R10975 iovss.n2473 iovss.n2398 4.49741
R10976 iovss.n2481 iovss.n2398 4.49741
R10977 iovss.n2423 iovss.n2398 4.49741
R10978 iovss.n2415 iovss.n2398 4.49741
R10979 iovss.n2497 iovss.n2398 4.49741
R10980 iovss.n2504 iovss.n2398 4.49741
R10981 iovss.n2455 iovss.n2399 4.49741
R10982 iovss.n2459 iovss.n2399 4.49741
R10983 iovss.n2450 iovss.n2399 4.49741
R10984 iovss.n2446 iovss.n2399 4.49741
R10985 iovss.n2442 iovss.n2399 4.49741
R10986 iovss.n2438 iovss.n2399 4.49741
R10987 iovss.n2471 iovss.n2399 4.49741
R10988 iovss.n2475 iovss.n2399 4.49741
R10989 iovss.n2479 iovss.n2399 4.49741
R10990 iovss.n2483 iovss.n2399 4.49741
R10991 iovss.n2425 iovss.n2399 4.49741
R10992 iovss.n2421 iovss.n2399 4.49741
R10993 iovss.n2417 iovss.n2399 4.49741
R10994 iovss.n2413 iovss.n2399 4.49741
R10995 iovss.n2495 iovss.n2399 4.49741
R10996 iovss.n2499 iovss.n2399 4.49741
R10997 iovss.n2506 iovss.n1444 4.49741
R10998 iovss.n2509 iovss.n2400 4.49741
R10999 iovss.n1991 iovss.n1990 4.49564
R11000 iovss.n1986 iovss.n1485 4.49564
R11001 iovss.n1991 iovss.n1989 4.49564
R11002 iovss.n1988 iovss.n1485 4.49564
R11003 iovss.n1542 iovss.n1535 4.49562
R11004 iovss.n1543 iovss.n1542 4.49562
R11005 iovss.n1547 iovss.n1534 4.49562
R11006 iovss.n1547 iovss.n1533 4.49562
R11007 iovss.n2932 iovss.n2931 4.49246
R11008 iovss.n2929 iovss.n2928 4.49246
R11009 iovss.n3071 iovss.n3070 4.49246
R11010 iovss.n3079 iovss.n2924 4.49246
R11011 iovss.n3070 iovss.n2937 4.49246
R11012 iovss.n3079 iovss.n2923 4.49246
R11013 iovss.n3070 iovss.n2938 4.49246
R11014 iovss.n3079 iovss.n2922 4.49246
R11015 iovss.n3070 iovss.n2939 4.49246
R11016 iovss.n3079 iovss.n2921 4.49246
R11017 iovss.n3070 iovss.n2940 4.49246
R11018 iovss.n3079 iovss.n2920 4.49246
R11019 iovss.n3070 iovss.n2941 4.49246
R11020 iovss.n3079 iovss.n2919 4.49246
R11021 iovss.n3070 iovss.n2942 4.49246
R11022 iovss.n3079 iovss.n2918 4.49246
R11023 iovss.n3070 iovss.n2943 4.49246
R11024 iovss.n3079 iovss.n2917 4.49246
R11025 iovss.n3070 iovss.n2944 4.49246
R11026 iovss.n3079 iovss.n2916 4.49246
R11027 iovss.n3070 iovss.n2945 4.49246
R11028 iovss.n3079 iovss.n2915 4.49246
R11029 iovss.n3070 iovss.n2946 4.49246
R11030 iovss.n3079 iovss.n2914 4.49246
R11031 iovss.n3070 iovss.n2947 4.49246
R11032 iovss.n3079 iovss.n2913 4.49246
R11033 iovss.n3070 iovss.n2948 4.49246
R11034 iovss.n3079 iovss.n2912 4.49246
R11035 iovss.n3070 iovss.n2949 4.49246
R11036 iovss.n3079 iovss.n2911 4.49246
R11037 iovss.n3070 iovss.n2950 4.49246
R11038 iovss.n3079 iovss.n2910 4.49246
R11039 iovss.n3070 iovss.n2951 4.49246
R11040 iovss.n3079 iovss.n2909 4.49246
R11041 iovss.n3070 iovss.n2952 4.49246
R11042 iovss.n3079 iovss.n2908 4.49246
R11043 iovss.n3070 iovss.n2953 4.49246
R11044 iovss.n3079 iovss.n2907 4.49246
R11045 iovss.n3070 iovss.n2954 4.49246
R11046 iovss.n3079 iovss.n2906 4.49246
R11047 iovss.n3070 iovss.n2955 4.49246
R11048 iovss.n3079 iovss.n2905 4.49246
R11049 iovss.n3070 iovss.n2956 4.49246
R11050 iovss.n3079 iovss.n2904 4.49246
R11051 iovss.n3070 iovss.n2957 4.49246
R11052 iovss.n3079 iovss.n2903 4.49246
R11053 iovss.n3070 iovss.n2958 4.49246
R11054 iovss.n3079 iovss.n2902 4.49246
R11055 iovss.n3070 iovss.n2927 4.49246
R11056 iovss.n1139 iovss.n1115 4.49246
R11057 iovss.n3095 iovss.n1109 4.49246
R11058 iovss.n3084 iovss.n1115 4.49246
R11059 iovss.n3098 iovss.n1142 4.49246
R11060 iovss.n1143 iovss.n1115 4.49246
R11061 iovss.n1145 iovss.n1115 4.49246
R11062 iovss.n1148 iovss.n1115 4.49246
R11063 iovss.n1151 iovss.n1115 4.49246
R11064 iovss.n1215 iovss.n1115 4.49246
R11065 iovss.n3098 iovss.n1131 4.49246
R11066 iovss.n1157 iovss.n1115 4.49246
R11067 iovss.n1159 iovss.n1115 4.49246
R11068 iovss.n3088 iovss.n1115 4.49246
R11069 iovss.n3098 iovss.n1162 4.49246
R11070 iovss.n1163 iovss.n1115 4.49246
R11071 iovss.n1165 iovss.n1115 4.49246
R11072 iovss.n1168 iovss.n1115 4.49246
R11073 iovss.n1171 iovss.n1115 4.49246
R11074 iovss.n1211 iovss.n1115 4.49246
R11075 iovss.n3098 iovss.n1123 4.49246
R11076 iovss.n1177 iovss.n1115 4.49246
R11077 iovss.n1179 iovss.n1115 4.49246
R11078 iovss.n3092 iovss.n1115 4.49246
R11079 iovss.n3098 iovss.n1182 4.49246
R11080 iovss.n1183 iovss.n1115 4.49246
R11081 iovss.n1185 iovss.n1115 4.49246
R11082 iovss.n1188 iovss.n1115 4.49246
R11083 iovss.n3099 iovss.n3098 4.49246
R11084 iovss.n3109 iovss.n988 4.49246
R11085 iovss.n1102 iovss.n1056 4.49246
R11086 iovss.n990 iovss.n962 4.49246
R11087 iovss.n1056 iovss.n1035 4.49246
R11088 iovss.n992 iovss.n962 4.49246
R11089 iovss.n1056 iovss.n1036 4.49246
R11090 iovss.n994 iovss.n962 4.49246
R11091 iovss.n1056 iovss.n1037 4.49246
R11092 iovss.n996 iovss.n962 4.49246
R11093 iovss.n1056 iovss.n1038 4.49246
R11094 iovss.n998 iovss.n962 4.49246
R11095 iovss.n1056 iovss.n1039 4.49246
R11096 iovss.n1000 iovss.n962 4.49246
R11097 iovss.n1056 iovss.n1040 4.49246
R11098 iovss.n1002 iovss.n962 4.49246
R11099 iovss.n1056 iovss.n1041 4.49246
R11100 iovss.n1004 iovss.n962 4.49246
R11101 iovss.n1056 iovss.n1042 4.49246
R11102 iovss.n1006 iovss.n962 4.49246
R11103 iovss.n1056 iovss.n1043 4.49246
R11104 iovss.n1008 iovss.n962 4.49246
R11105 iovss.n1056 iovss.n1044 4.49246
R11106 iovss.n1010 iovss.n962 4.49246
R11107 iovss.n1056 iovss.n1045 4.49246
R11108 iovss.n1012 iovss.n962 4.49246
R11109 iovss.n1056 iovss.n1046 4.49246
R11110 iovss.n1014 iovss.n962 4.49246
R11111 iovss.n1056 iovss.n1047 4.49246
R11112 iovss.n1016 iovss.n962 4.49246
R11113 iovss.n1056 iovss.n1048 4.49246
R11114 iovss.n1018 iovss.n962 4.49246
R11115 iovss.n1056 iovss.n1049 4.49246
R11116 iovss.n1020 iovss.n962 4.49246
R11117 iovss.n1056 iovss.n1050 4.49246
R11118 iovss.n1022 iovss.n962 4.49246
R11119 iovss.n1056 iovss.n1051 4.49246
R11120 iovss.n1024 iovss.n962 4.49246
R11121 iovss.n1056 iovss.n1052 4.49246
R11122 iovss.n1026 iovss.n962 4.49246
R11123 iovss.n1056 iovss.n1053 4.49246
R11124 iovss.n1028 iovss.n962 4.49246
R11125 iovss.n1056 iovss.n1054 4.49246
R11126 iovss.n1030 iovss.n962 4.49246
R11127 iovss.n1056 iovss.n1055 4.49246
R11128 iovss.n1032 iovss.n962 4.49246
R11129 iovss.n1056 iovss.n963 4.49246
R11130 iovss.n3111 iovss.n962 4.49246
R11131 iovss.n2900 iovss.n1226 4.49246
R11132 iovss.n2886 iovss.n2790 4.49246
R11133 iovss.n2900 iovss.n1227 4.49246
R11134 iovss.n2886 iovss.n2795 4.49246
R11135 iovss.n2900 iovss.n1228 4.49246
R11136 iovss.n2886 iovss.n2800 4.49246
R11137 iovss.n2900 iovss.n1229 4.49246
R11138 iovss.n2886 iovss.n2805 4.49246
R11139 iovss.n2900 iovss.n1230 4.49246
R11140 iovss.n2886 iovss.n2810 4.49246
R11141 iovss.n2900 iovss.n1231 4.49246
R11142 iovss.n2886 iovss.n2815 4.49246
R11143 iovss.n2900 iovss.n1232 4.49246
R11144 iovss.n2886 iovss.n2820 4.49246
R11145 iovss.n2900 iovss.n1233 4.49246
R11146 iovss.n2886 iovss.n2825 4.49246
R11147 iovss.n2900 iovss.n1234 4.49246
R11148 iovss.n2886 iovss.n2830 4.49246
R11149 iovss.n2900 iovss.n1235 4.49246
R11150 iovss.n2886 iovss.n2835 4.49246
R11151 iovss.n2900 iovss.n1236 4.49246
R11152 iovss.n2886 iovss.n2840 4.49246
R11153 iovss.n2900 iovss.n1237 4.49246
R11154 iovss.n2886 iovss.n2845 4.49246
R11155 iovss.n2900 iovss.n1238 4.49246
R11156 iovss.n2886 iovss.n2850 4.49246
R11157 iovss.n2900 iovss.n1239 4.49246
R11158 iovss.n2886 iovss.n2855 4.49246
R11159 iovss.n2900 iovss.n1240 4.49246
R11160 iovss.n2886 iovss.n2860 4.49246
R11161 iovss.n2900 iovss.n1241 4.49246
R11162 iovss.n2886 iovss.n2865 4.49246
R11163 iovss.n2900 iovss.n1242 4.49246
R11164 iovss.n2886 iovss.n2870 4.49246
R11165 iovss.n2900 iovss.n1243 4.49246
R11166 iovss.n2886 iovss.n2875 4.49246
R11167 iovss.n2900 iovss.n1244 4.49246
R11168 iovss.n2886 iovss.n2880 4.49246
R11169 iovss.n2900 iovss.n1245 4.49246
R11170 iovss.n2886 iovss.n2885 4.49246
R11171 iovss.n2900 iovss.n1246 4.49246
R11172 iovss.n2888 iovss.n2886 4.49246
R11173 iovss.n2886 iovss.n1247 4.49246
R11174 iovss.n2898 iovss.n1219 4.49246
R11175 iovss.n2751 iovss.n1409 4.49246
R11176 iovss.n2647 iovss.n2602 4.49246
R11177 iovss.n2751 iovss.n2730 4.49246
R11178 iovss.n2650 iovss.n2602 4.49246
R11179 iovss.n2751 iovss.n2731 4.49246
R11180 iovss.n2653 iovss.n2602 4.49246
R11181 iovss.n2751 iovss.n2732 4.49246
R11182 iovss.n2656 iovss.n2602 4.49246
R11183 iovss.n2751 iovss.n2733 4.49246
R11184 iovss.n2659 iovss.n2602 4.49246
R11185 iovss.n2751 iovss.n2734 4.49246
R11186 iovss.n2662 iovss.n2602 4.49246
R11187 iovss.n2751 iovss.n2735 4.49246
R11188 iovss.n2665 iovss.n2602 4.49246
R11189 iovss.n2751 iovss.n2736 4.49246
R11190 iovss.n2668 iovss.n2602 4.49246
R11191 iovss.n2751 iovss.n2737 4.49246
R11192 iovss.n2671 iovss.n2602 4.49246
R11193 iovss.n2751 iovss.n2738 4.49246
R11194 iovss.n2674 iovss.n2602 4.49246
R11195 iovss.n2751 iovss.n2739 4.49246
R11196 iovss.n2677 iovss.n2602 4.49246
R11197 iovss.n2751 iovss.n2740 4.49246
R11198 iovss.n2680 iovss.n2602 4.49246
R11199 iovss.n2751 iovss.n2741 4.49246
R11200 iovss.n2683 iovss.n2602 4.49246
R11201 iovss.n2751 iovss.n2742 4.49246
R11202 iovss.n2686 iovss.n2602 4.49246
R11203 iovss.n2751 iovss.n2743 4.49246
R11204 iovss.n2689 iovss.n2602 4.49246
R11205 iovss.n2751 iovss.n2744 4.49246
R11206 iovss.n2692 iovss.n2602 4.49246
R11207 iovss.n2751 iovss.n2745 4.49246
R11208 iovss.n2695 iovss.n2602 4.49246
R11209 iovss.n2751 iovss.n2746 4.49246
R11210 iovss.n2698 iovss.n2602 4.49246
R11211 iovss.n2751 iovss.n2747 4.49246
R11212 iovss.n2701 iovss.n2602 4.49246
R11213 iovss.n2751 iovss.n2748 4.49246
R11214 iovss.n2704 iovss.n2602 4.49246
R11215 iovss.n2751 iovss.n2749 4.49246
R11216 iovss.n2707 iovss.n2602 4.49246
R11217 iovss.n2751 iovss.n2750 4.49246
R11218 iovss.n2710 iovss.n2602 4.49246
R11219 iovss.n2760 iovss.n1344 4.49246
R11220 iovss.n1380 iovss.n1341 4.49246
R11221 iovss.n1345 iovss.n1340 4.49246
R11222 iovss.n1348 iovss.n1341 4.49246
R11223 iovss.n1347 iovss.n1340 4.49246
R11224 iovss.n1341 iovss.n1338 4.49246
R11225 iovss.n2768 iovss.n1312 4.49246
R11226 iovss.n2764 iovss.n1309 4.49246
R11227 iovss.n2771 iovss.n1312 4.49246
R11228 iovss.n2766 iovss.n1309 4.49246
R11229 iovss.n2775 iovss.n1312 4.49246
R11230 iovss.n1313 iovss.n1309 4.49246
R11231 iovss.n893 iovss.n886 4.49246
R11232 iovss.n3144 iovss.n3139 4.49246
R11233 iovss.n895 iovss.n886 4.49246
R11234 iovss.n3144 iovss.n3140 4.49246
R11235 iovss.n897 iovss.n886 4.49246
R11236 iovss.n3144 iovss.n3141 4.49246
R11237 iovss.n899 iovss.n886 4.49246
R11238 iovss.n3144 iovss.n3142 4.49246
R11239 iovss.n901 iovss.n886 4.49246
R11240 iovss.n3144 iovss.n3143 4.49246
R11241 iovss.n903 iovss.n886 4.49246
R11242 iovss.n1198 iovss.n1196 4.49246
R11243 iovss.n916 iovss.n907 4.49246
R11244 iovss.n1198 iovss.n1197 4.49246
R11245 iovss.n921 iovss.n907 4.49246
R11246 iovss.n1198 iovss.n1195 4.49246
R11247 iovss.n1198 iovss.n926 4.49246
R11248 iovss.n925 iovss.n907 4.49246
R11249 iovss.n1198 iovss.n906 4.49246
R11250 iovss.n939 iovss.n930 4.49246
R11251 iovss.n949 iovss.n946 4.49246
R11252 iovss.n941 iovss.n930 4.49246
R11253 iovss.n949 iovss.n947 4.49246
R11254 iovss.n943 iovss.n930 4.49246
R11255 iovss.n949 iovss.n948 4.49246
R11256 iovss.n951 iovss.n930 4.49246
R11257 iovss.n950 iovss.n949 4.49246
R11258 iovss.n930 iovss.n929 4.49246
R11259 iovss.n949 iovss.n928 4.49246
R11260 iovss.n931 iovss.n930 4.49246
R11261 iovss.n3103 iovss.t3 3.07412
R11262 iovss.n1110 iovss.t1 3.07412
R11263 iovss.n2761 iovss.n1339 3.02695
R11264 iovss.n2765 iovss.n1277 3.02695
R11265 iovss.n578 iovss.n577 3.023
R11266 iovss.n3466 iovss.n3464 3.0115
R11267 iovss.n1216 iovss.n904 3.00792
R11268 iovss.n911 iovss.n904 3.0079
R11269 iovss.n3093 iovss.n904 3.0079
R11270 iovss.n1212 iovss.n904 3.00782
R11271 iovss.n3089 iovss.n904 3.00769
R11272 iovss.n3085 iovss.n904 3.00728
R11273 iovss.n3135 iovss.n3134 3.00565
R11274 iovss.n1138 iovss.n1137 3.00498
R11275 iovss.n915 iovss.n904 3.00422
R11276 iovss.n3113 iovss.n960 3.0005
R11277 iovss.n959 iovss.n957 3.0005
R11278 iovss.n3117 iovss.n956 3.0005
R11279 iovss.n3118 iovss.n955 3.0005
R11280 iovss.n3119 iovss.n954 3.0005
R11281 iovss.n1107 iovss.n1106 3.0005
R11282 iovss.n3132 iovss.n3131 3.0005
R11283 iovss.n952 iovss.n934 3.0005
R11284 iovss.n3129 iovss.n3128 3.0005
R11285 iovss.n3127 iovss.n935 3.0005
R11286 iovss.n3126 iovss.n944 3.0005
R11287 iovss.n3125 iovss.n936 3.0005
R11288 iovss.n3124 iovss.n942 3.0005
R11289 iovss.n3123 iovss.n937 3.0005
R11290 iovss.n3122 iovss.n940 3.0005
R11291 iovss.n3121 iovss.n938 3.0005
R11292 iovss.n3120 iovss.n3119 3.0005
R11293 iovss.n3118 iovss.n953 3.0005
R11294 iovss.n3117 iovss.n3116 3.0005
R11295 iovss.n3115 iovss.n957 3.0005
R11296 iovss.n3114 iovss.n3113 3.0005
R11297 iovss.n3112 iovss.n958 3.0005
R11298 iovss.n3110 iovss.n964 3.0005
R11299 iovss.n1058 iovss.n1033 3.0005
R11300 iovss.n1059 iovss.n966 3.0005
R11301 iovss.n1060 iovss.n1031 3.0005
R11302 iovss.n1061 iovss.n967 3.0005
R11303 iovss.n1062 iovss.n1029 3.0005
R11304 iovss.n1063 iovss.n968 3.0005
R11305 iovss.n1064 iovss.n1027 3.0005
R11306 iovss.n1065 iovss.n969 3.0005
R11307 iovss.n1066 iovss.n1025 3.0005
R11308 iovss.n1067 iovss.n970 3.0005
R11309 iovss.n1068 iovss.n1023 3.0005
R11310 iovss.n1069 iovss.n971 3.0005
R11311 iovss.n1070 iovss.n1021 3.0005
R11312 iovss.n1071 iovss.n972 3.0005
R11313 iovss.n1072 iovss.n1019 3.0005
R11314 iovss.n1073 iovss.n973 3.0005
R11315 iovss.n1074 iovss.n1017 3.0005
R11316 iovss.n1075 iovss.n974 3.0005
R11317 iovss.n1076 iovss.n1015 3.0005
R11318 iovss.n1077 iovss.n975 3.0005
R11319 iovss.n1078 iovss.n1013 3.0005
R11320 iovss.n1079 iovss.n976 3.0005
R11321 iovss.n1080 iovss.n1011 3.0005
R11322 iovss.n1081 iovss.n977 3.0005
R11323 iovss.n1082 iovss.n1009 3.0005
R11324 iovss.n1083 iovss.n978 3.0005
R11325 iovss.n1084 iovss.n1007 3.0005
R11326 iovss.n1085 iovss.n979 3.0005
R11327 iovss.n1086 iovss.n1005 3.0005
R11328 iovss.n1087 iovss.n980 3.0005
R11329 iovss.n1088 iovss.n1003 3.0005
R11330 iovss.n1089 iovss.n981 3.0005
R11331 iovss.n1090 iovss.n1001 3.0005
R11332 iovss.n1091 iovss.n982 3.0005
R11333 iovss.n1092 iovss.n999 3.0005
R11334 iovss.n1093 iovss.n983 3.0005
R11335 iovss.n1094 iovss.n997 3.0005
R11336 iovss.n1095 iovss.n984 3.0005
R11337 iovss.n1096 iovss.n995 3.0005
R11338 iovss.n1097 iovss.n985 3.0005
R11339 iovss.n1098 iovss.n993 3.0005
R11340 iovss.n1099 iovss.n986 3.0005
R11341 iovss.n1100 iovss.n991 3.0005
R11342 iovss.n1101 iovss.n987 3.0005
R11343 iovss.n1104 iovss.n1103 3.0005
R11344 iovss.n3138 iovss.n905 3.0005
R11345 iovss.n933 iovss.n932 3.0005
R11346 iovss.n3138 iovss.n3137 3.0005
R11347 iovss.n932 iovss.n908 3.0005
R11348 iovss.n1207 iovss.n1206 3.0005
R11349 iovss.n1205 iovss.n1204 3.0005
R11350 iovss.n1203 iovss.n1192 3.0005
R11351 iovss.n1201 iovss.n1200 3.0005
R11352 iovss.n1199 iovss.n1194 3.0005
R11353 iovss.n3075 iovss.n2925 3.0005
R11354 iovss.n2966 iovss.n889 3.0005
R11355 iovss.n2967 iovss.n898 3.0005
R11356 iovss.n2968 iovss.n890 3.0005
R11357 iovss.n2969 iovss.n896 3.0005
R11358 iovss.n2970 iovss.n891 3.0005
R11359 iovss.n2971 iovss.n894 3.0005
R11360 iovss.n2972 iovss.n892 3.0005
R11361 iovss.n2973 iovss.n2963 3.0005
R11362 iovss.n2975 iovss.n2974 3.0005
R11363 iovss.n2961 iovss.n2960 3.0005
R11364 iovss.n2980 iovss.n2979 3.0005
R11365 iovss.n2981 iovss.n2959 3.0005
R11366 iovss.n3069 iovss.n3068 3.0005
R11367 iovss.n3067 iovss.n3066 3.0005
R11368 iovss.n3065 iovss.n3064 3.0005
R11369 iovss.n3063 iovss.n3062 3.0005
R11370 iovss.n3061 iovss.n3060 3.0005
R11371 iovss.n3059 iovss.n3058 3.0005
R11372 iovss.n3057 iovss.n3056 3.0005
R11373 iovss.n3055 iovss.n3054 3.0005
R11374 iovss.n3053 iovss.n3052 3.0005
R11375 iovss.n3051 iovss.n3050 3.0005
R11376 iovss.n3049 iovss.n3048 3.0005
R11377 iovss.n3047 iovss.n3046 3.0005
R11378 iovss.n3045 iovss.n3044 3.0005
R11379 iovss.n3043 iovss.n3042 3.0005
R11380 iovss.n3041 iovss.n3040 3.0005
R11381 iovss.n3039 iovss.n3038 3.0005
R11382 iovss.n3037 iovss.n3036 3.0005
R11383 iovss.n3035 iovss.n3034 3.0005
R11384 iovss.n3033 iovss.n3032 3.0005
R11385 iovss.n3031 iovss.n3030 3.0005
R11386 iovss.n3029 iovss.n3028 3.0005
R11387 iovss.n3027 iovss.n3026 3.0005
R11388 iovss.n3025 iovss.n3024 3.0005
R11389 iovss.n3023 iovss.n3022 3.0005
R11390 iovss.n3021 iovss.n3020 3.0005
R11391 iovss.n3019 iovss.n3018 3.0005
R11392 iovss.n3017 iovss.n3016 3.0005
R11393 iovss.n3015 iovss.n3014 3.0005
R11394 iovss.n3013 iovss.n3012 3.0005
R11395 iovss.n3011 iovss.n3010 3.0005
R11396 iovss.n3009 iovss.n3008 3.0005
R11397 iovss.n3007 iovss.n3006 3.0005
R11398 iovss.n3005 iovss.n3004 3.0005
R11399 iovss.n3003 iovss.n3002 3.0005
R11400 iovss.n3001 iovss.n3000 3.0005
R11401 iovss.n2999 iovss.n2998 3.0005
R11402 iovss.n2997 iovss.n2996 3.0005
R11403 iovss.n2995 iovss.n2994 3.0005
R11404 iovss.n2993 iovss.n2992 3.0005
R11405 iovss.n2991 iovss.n2990 3.0005
R11406 iovss.n2989 iovss.n2988 3.0005
R11407 iovss.n2987 iovss.n2986 3.0005
R11408 iovss.n2985 iovss.n2984 3.0005
R11409 iovss.n2983 iovss.n2982 3.0005
R11410 iovss.n2936 iovss.n2933 3.0005
R11411 iovss.n3073 iovss.n3072 3.0005
R11412 iovss.n3074 iovss.n2926 3.0005
R11413 iovss.n927 iovss.n902 3.0005
R11414 iovss.n3145 iovss.n3138 3.0005
R11415 iovss.n932 iovss.n887 3.0005
R11416 iovss.n2964 iovss.n888 3.0005
R11417 iovss.n2965 iovss.n900 3.0005
R11418 iovss.n2959 iovss.n2934 3.0005
R11419 iovss.n2979 iovss.n2978 3.0005
R11420 iovss.n2977 iovss.n2961 3.0005
R11421 iovss.n2976 iovss.n2975 3.0005
R11422 iovss.n2963 iovss.n2962 3.0005
R11423 iovss.n579 iovss.n576 3.0005
R11424 iovss.n581 iovss.n573 3.0005
R11425 iovss.n584 iovss.n583 3.0005
R11426 iovss.n569 iovss.n568 3.0005
R11427 iovss.n594 iovss.n592 3.0005
R11428 iovss.n597 iovss.n596 3.0005
R11429 iovss.n598 iovss.n559 3.0005
R11430 iovss.n607 iovss.n606 3.0005
R11431 iovss.n562 iovss.n488 3.0005
R11432 iovss.n3261 iovss.n486 3.0005
R11433 iovss.n3263 iovss.n3262 3.0005
R11434 iovss.n482 iovss.n481 3.0005
R11435 iovss.n3274 iovss.n3272 3.0005
R11436 iovss.n3276 iovss.n479 3.0005
R11437 iovss.n3279 iovss.n3278 3.0005
R11438 iovss.n475 iovss.n474 3.0005
R11439 iovss.n3289 iovss.n3287 3.0005
R11440 iovss.n3292 iovss.n3291 3.0005
R11441 iovss.n3294 iovss.n453 3.0005
R11442 iovss.n3337 iovss.n454 3.0005
R11443 iovss.n3336 iovss.n455 3.0005
R11444 iovss.n3332 iovss.n456 3.0005
R11445 iovss.n3331 iovss.n457 3.0005
R11446 iovss.n3329 iovss.n458 3.0005
R11447 iovss.n3327 iovss.n459 3.0005
R11448 iovss.n3326 iovss.n460 3.0005
R11449 iovss.n3324 iovss.n461 3.0005
R11450 iovss.n3322 iovss.n3320 3.0005
R11451 iovss.n463 iovss.n77 3.0005
R11452 iovss.n3439 iovss.n3438 3.0005
R11453 iovss.n3440 iovss.n69 3.0005
R11454 iovss.n3450 iovss.n3449 3.0005
R11455 iovss.n71 iovss.n67 3.0005
R11456 iovss.n3455 iovss.n3454 3.0005
R11457 iovss.n3457 iovss.n59 3.0005
R11458 iovss.n3469 iovss.n60 3.0005
R11459 iovss.n3468 iovss.n61 3.0005
R11460 iovss.n3466 iovss.n3465 3.0005
R11461 iovss.n3468 iovss.n3467 3.0005
R11462 iovss.n3470 iovss.n3469 3.0005
R11463 iovss.n59 iovss.n58 3.0005
R11464 iovss.n3454 iovss.n3453 3.0005
R11465 iovss.n3452 iovss.n67 3.0005
R11466 iovss.n3451 iovss.n3450 3.0005
R11467 iovss.n94 iovss.n69 3.0005
R11468 iovss.n3438 iovss.n3437 3.0005
R11469 iovss.n144 iovss.n77 3.0005
R11470 iovss.n3322 iovss.n3321 3.0005
R11471 iovss.n3324 iovss.n3323 3.0005
R11472 iovss.n3326 iovss.n3325 3.0005
R11473 iovss.n3327 iovss.n113 3.0005
R11474 iovss.n3329 iovss.n3328 3.0005
R11475 iovss.n3331 iovss.n3330 3.0005
R11476 iovss.n3334 iovss.n3332 3.0005
R11477 iovss.n3336 iovss.n3335 3.0005
R11478 iovss.n3338 iovss.n3337 3.0005
R11479 iovss.n453 iovss.n452 3.0005
R11480 iovss.n3291 iovss.n3290 3.0005
R11481 iovss.n3289 iovss.n3288 3.0005
R11482 iovss.n474 iovss.n473 3.0005
R11483 iovss.n3278 iovss.n3277 3.0005
R11484 iovss.n3276 iovss.n3275 3.0005
R11485 iovss.n3274 iovss.n3273 3.0005
R11486 iovss.n481 iovss.n388 3.0005
R11487 iovss.n3262 iovss.n380 3.0005
R11488 iovss.n3261 iovss.n3260 3.0005
R11489 iovss.n612 iovss.n488 3.0005
R11490 iovss.n608 iovss.n607 3.0005
R11491 iovss.n559 iovss.n558 3.0005
R11492 iovss.n596 iovss.n595 3.0005
R11493 iovss.n594 iovss.n593 3.0005
R11494 iovss.n568 iovss.n567 3.0005
R11495 iovss.n583 iovss.n582 3.0005
R11496 iovss.n581 iovss.n580 3.0005
R11497 iovss.n2899 iovss.n1248 3.0005
R11498 iovss.n2893 iovss.n2892 3.0005
R11499 iovss.n2890 iovss.n2889 3.0005
R11500 iovss.n2887 iovss.n1304 3.0005
R11501 iovss.n2882 iovss.n2881 3.0005
R11502 iovss.n2884 iovss.n2883 3.0005
R11503 iovss.n2877 iovss.n2876 3.0005
R11504 iovss.n2879 iovss.n2878 3.0005
R11505 iovss.n2872 iovss.n2871 3.0005
R11506 iovss.n2874 iovss.n2873 3.0005
R11507 iovss.n2867 iovss.n2866 3.0005
R11508 iovss.n2869 iovss.n2868 3.0005
R11509 iovss.n2862 iovss.n2861 3.0005
R11510 iovss.n2864 iovss.n2863 3.0005
R11511 iovss.n2857 iovss.n2856 3.0005
R11512 iovss.n2859 iovss.n2858 3.0005
R11513 iovss.n2852 iovss.n2851 3.0005
R11514 iovss.n2854 iovss.n2853 3.0005
R11515 iovss.n2847 iovss.n2846 3.0005
R11516 iovss.n2849 iovss.n2848 3.0005
R11517 iovss.n2842 iovss.n2841 3.0005
R11518 iovss.n2844 iovss.n2843 3.0005
R11519 iovss.n2837 iovss.n2836 3.0005
R11520 iovss.n2839 iovss.n2838 3.0005
R11521 iovss.n2832 iovss.n2831 3.0005
R11522 iovss.n2834 iovss.n2833 3.0005
R11523 iovss.n2827 iovss.n2826 3.0005
R11524 iovss.n2829 iovss.n2828 3.0005
R11525 iovss.n2822 iovss.n2821 3.0005
R11526 iovss.n2824 iovss.n2823 3.0005
R11527 iovss.n2817 iovss.n2816 3.0005
R11528 iovss.n2819 iovss.n2818 3.0005
R11529 iovss.n2812 iovss.n2811 3.0005
R11530 iovss.n2814 iovss.n2813 3.0005
R11531 iovss.n2807 iovss.n2806 3.0005
R11532 iovss.n2809 iovss.n2808 3.0005
R11533 iovss.n2802 iovss.n2801 3.0005
R11534 iovss.n2804 iovss.n2803 3.0005
R11535 iovss.n2797 iovss.n2796 3.0005
R11536 iovss.n2799 iovss.n2798 3.0005
R11537 iovss.n2792 iovss.n2791 3.0005
R11538 iovss.n2794 iovss.n2793 3.0005
R11539 iovss.n2789 iovss.n2788 3.0005
R11540 iovss.n1284 iovss.n1225 3.0005
R11541 iovss.n2786 iovss.n2785 3.0005
R11542 iovss.n2784 iovss.n2783 3.0005
R11543 iovss.n2782 iovss.n1308 3.0005
R11544 iovss.n1307 iovss.n1306 3.0005
R11545 iovss.n2778 iovss.n2777 3.0005
R11546 iovss.n2776 iovss.n1311 3.0005
R11547 iovss.n2774 iovss.n1314 3.0005
R11548 iovss.n2772 iovss.n2770 3.0005
R11549 iovss.n1316 iovss.n1315 3.0005
R11550 iovss.n2769 iovss.n2767 3.0005
R11551 iovss.n1318 iovss.n1317 3.0005
R11552 iovss.n2779 iovss.n2778 3.0005
R11553 iovss.n2780 iovss.n1307 3.0005
R11554 iovss.n2782 iovss.n2781 3.0005
R11555 iovss.n2784 iovss.n1305 3.0005
R11556 iovss.n2787 iovss.n2786 3.0005
R11557 iovss.n2897 iovss.n2896 3.0005
R11558 iovss.n2645 iovss.n1408 3.0005
R11559 iovss.n2648 iovss.n2646 3.0005
R11560 iovss.n2644 iovss.n2643 3.0005
R11561 iovss.n2651 iovss.n2649 3.0005
R11562 iovss.n2642 iovss.n2641 3.0005
R11563 iovss.n2654 iovss.n2652 3.0005
R11564 iovss.n2640 iovss.n2639 3.0005
R11565 iovss.n2657 iovss.n2655 3.0005
R11566 iovss.n2638 iovss.n2637 3.0005
R11567 iovss.n2660 iovss.n2658 3.0005
R11568 iovss.n2636 iovss.n2635 3.0005
R11569 iovss.n2663 iovss.n2661 3.0005
R11570 iovss.n2634 iovss.n2633 3.0005
R11571 iovss.n2666 iovss.n2664 3.0005
R11572 iovss.n2632 iovss.n2631 3.0005
R11573 iovss.n2669 iovss.n2667 3.0005
R11574 iovss.n2630 iovss.n2629 3.0005
R11575 iovss.n2672 iovss.n2670 3.0005
R11576 iovss.n2628 iovss.n2627 3.0005
R11577 iovss.n2675 iovss.n2673 3.0005
R11578 iovss.n2626 iovss.n2625 3.0005
R11579 iovss.n2678 iovss.n2676 3.0005
R11580 iovss.n2624 iovss.n2623 3.0005
R11581 iovss.n2681 iovss.n2679 3.0005
R11582 iovss.n2622 iovss.n2621 3.0005
R11583 iovss.n2684 iovss.n2682 3.0005
R11584 iovss.n2620 iovss.n2619 3.0005
R11585 iovss.n2687 iovss.n2685 3.0005
R11586 iovss.n2618 iovss.n2617 3.0005
R11587 iovss.n2690 iovss.n2688 3.0005
R11588 iovss.n2616 iovss.n2615 3.0005
R11589 iovss.n2693 iovss.n2691 3.0005
R11590 iovss.n2614 iovss.n2613 3.0005
R11591 iovss.n2696 iovss.n2694 3.0005
R11592 iovss.n2612 iovss.n2611 3.0005
R11593 iovss.n2699 iovss.n2697 3.0005
R11594 iovss.n2610 iovss.n2609 3.0005
R11595 iovss.n2702 iovss.n2700 3.0005
R11596 iovss.n2608 iovss.n2607 3.0005
R11597 iovss.n2705 iovss.n2703 3.0005
R11598 iovss.n2606 iovss.n2605 3.0005
R11599 iovss.n2708 iovss.n2706 3.0005
R11600 iovss.n2604 iovss.n2603 3.0005
R11601 iovss.n2711 iovss.n2709 3.0005
R11602 iovss.n2728 iovss.n2727 3.0005
R11603 iovss.n2726 iovss.n2725 3.0005
R11604 iovss.n2724 iovss.n2715 3.0005
R11605 iovss.n2714 iovss.n2713 3.0005
R11606 iovss.n2720 iovss.n2719 3.0005
R11607 iovss.n2718 iovss.n2717 3.0005
R11608 iovss.n1382 iovss.n1381 3.0005
R11609 iovss.n1378 iovss.n1346 3.0005
R11610 iovss.n1351 iovss.n1343 3.0005
R11611 iovss.n2759 iovss.n2758 3.0005
R11612 iovss.n1349 iovss.n1342 3.0005
R11613 iovss.n2755 iovss.n2754 3.0005
R11614 iovss.n2729 iovss.n2728 3.0005
R11615 iovss.n2726 iovss.n2712 3.0005
R11616 iovss.n2724 iovss.n2723 3.0005
R11617 iovss.n2722 iovss.n2714 3.0005
R11618 iovss.n2721 iovss.n2720 3.0005
R11619 iovss.t2 iovss.n1364 2.82732
R11620 iovss.t0 iovss.n1262 2.82732
R11621 iovss.t2 iovss.n1339 2.82704
R11622 iovss.t0 iovss.n1277 2.82704
R11623 iovss.t2 iovss.n1377 2.82693
R11624 iovss.t2 iovss.n1383 2.82693
R11625 iovss.t2 iovss.n1375 2.82693
R11626 iovss.t2 iovss.n1385 2.82693
R11627 iovss.t2 iovss.n1387 2.82693
R11628 iovss.t2 iovss.n1372 2.82693
R11629 iovss.t2 iovss.n1389 2.82693
R11630 iovss.t2 iovss.n1370 2.82693
R11631 iovss.t2 iovss.n1368 2.82693
R11632 iovss.t2 iovss.n1392 2.82693
R11633 iovss.t2 iovss.n1366 2.82693
R11634 iovss.t2 iovss.n1395 2.82693
R11635 iovss.t2 iovss.n1362 2.82693
R11636 iovss.t2 iovss.n1397 2.82693
R11637 iovss.t2 iovss.n1399 2.82693
R11638 iovss.t2 iovss.n1359 2.82693
R11639 iovss.t2 iovss.n1401 2.82693
R11640 iovss.t2 iovss.n1357 2.82693
R11641 iovss.t2 iovss.n1355 2.82693
R11642 iovss.t2 iovss.n1404 2.82693
R11643 iovss.t2 iovss.n1353 2.82693
R11644 iovss.t2 iovss.n1406 2.82693
R11645 iovss.t2 iovss.n2756 2.82693
R11646 iovss.t0 iovss.n1275 2.82693
R11647 iovss.t0 iovss.n1280 2.82693
R11648 iovss.t0 iovss.n1273 2.82693
R11649 iovss.t0 iovss.n1282 2.82693
R11650 iovss.t0 iovss.n1285 2.82693
R11651 iovss.t0 iovss.n1270 2.82693
R11652 iovss.t0 iovss.n1287 2.82693
R11653 iovss.t0 iovss.n1268 2.82693
R11654 iovss.t0 iovss.n1266 2.82693
R11655 iovss.t0 iovss.n1290 2.82693
R11656 iovss.t0 iovss.n1264 2.82693
R11657 iovss.t0 iovss.n1293 2.82693
R11658 iovss.t0 iovss.n1260 2.82693
R11659 iovss.t0 iovss.n1295 2.82693
R11660 iovss.t0 iovss.n1297 2.82693
R11661 iovss.t0 iovss.n1257 2.82693
R11662 iovss.t0 iovss.n1299 2.82693
R11663 iovss.t0 iovss.n1255 2.82693
R11664 iovss.t0 iovss.n1253 2.82693
R11665 iovss.t0 iovss.n1302 2.82693
R11666 iovss.t0 iovss.n1251 2.82693
R11667 iovss.t0 iovss.n2891 2.82693
R11668 iovss.n2895 iovss.t0 2.82693
R11669 iovss.n2038 iovss.n2034 2.20699
R11670 iovss.n2593 iovss.n1428 2.20699
R11671 iovss.n2595 iovss.n2594 2.2005
R11672 iovss.n1429 iovss.n1427 2.2005
R11673 iovss.n2590 iovss.n2589 2.2005
R11674 iovss.n1432 iovss.n1431 2.2005
R11675 iovss.n2436 iovss.n2435 2.2005
R11676 iovss.n2464 iovss.n2463 2.2005
R11677 iovss.n2465 iovss.n2429 2.2005
R11678 iovss.n2467 iovss.n2466 2.2005
R11679 iovss.n2411 iovss.n2410 2.2005
R11680 iovss.n2488 iovss.n2487 2.2005
R11681 iovss.n2489 iovss.n2405 2.2005
R11682 iovss.n2491 iovss.n2490 2.2005
R11683 iovss.n1530 iovss.n1529 2.2005
R11684 iovss.n2514 iovss.n2513 2.2005
R11685 iovss.n2515 iovss.n1524 2.2005
R11686 iovss.n2517 iovss.n2516 2.2005
R11687 iovss.n1522 iovss.n1521 2.2005
R11688 iovss.n2524 iovss.n2523 2.2005
R11689 iovss.n2525 iovss.n1516 2.2005
R11690 iovss.n2527 iovss.n2526 2.2005
R11691 iovss.n1513 iovss.n1512 2.2005
R11692 iovss.n2535 iovss.n2534 2.2005
R11693 iovss.n2536 iovss.n1507 2.2005
R11694 iovss.n2538 iovss.n2537 2.2005
R11695 iovss.n1508 iovss.n1506 2.2005
R11696 iovss.n2053 iovss.n2052 2.2005
R11697 iovss.n2059 iovss.n2058 2.2005
R11698 iovss.n2060 iovss.n2045 2.2005
R11699 iovss.n2062 iovss.n2061 2.2005
R11700 iovss.n2042 iovss.n2041 2.2005
R11701 iovss.n2070 iovss.n2069 2.2005
R11702 iovss.n2071 iovss.n2037 2.2005
R11703 iovss.n2073 iovss.n2072 2.2005
R11704 iovss.n2762 iovss.n1320 1.67082
R11705 iovss.n2763 iovss.n1319 1.67082
R11706 iovss.n578 iovss.n537 1.51387
R11707 iovss.n1416 iovss.n1249 1.5005
R11708 iovss.n1424 iovss.n1423 1.5005
R11709 iovss.n1422 iovss.n1415 1.5005
R11710 iovss.n1421 iovss.n1420 1.5005
R11711 iovss.n1419 iovss.n1418 1.5005
R11712 iovss.n1417 iovss.n1413 1.5005
R11713 iovss.n2598 iovss.n1411 1.5005
R11714 iovss.n2600 iovss.n2599 1.5005
R11715 iovss.n1412 iovss.n1410 1.5005
R11716 iovss.n2579 iovss.n2578 1.5005
R11717 iovss.n2581 iovss.n2577 1.5005
R11718 iovss.n2583 iovss.n2582 1.5005
R11719 iovss.n2584 iovss.n1435 1.5005
R11720 iovss.n2586 iovss.n2585 1.5005
R11721 iovss.n2576 iovss.n1434 1.5005
R11722 iovss.n2575 iovss.n2574 1.5005
R11723 iovss.n2573 iovss.n1436 1.5005
R11724 iovss.n2572 iovss.n2571 1.5005
R11725 iovss.n2570 iovss.n2569 1.5005
R11726 iovss.n2568 iovss.n1438 1.5005
R11727 iovss.n2567 iovss.n2566 1.5005
R11728 iovss.n2565 iovss.n1439 1.5005
R11729 iovss.n1193 iovss.n904 1.49548
R11730 iovss.n1202 iovss.n904 1.49532
R11731 iovss.n923 iovss.n904 1.49504
R11732 iovss.n1176 iovss.n904 1.49504
R11733 iovss.n1169 iovss.n904 1.49504
R11734 iovss.n1140 iovss.n904 1.49504
R11735 iovss.n1189 iovss.n904 1.49502
R11736 iovss.n1156 iovss.n904 1.49502
R11737 iovss.n1152 iovss.n904 1.49502
R11738 iovss.n1186 iovss.n904 1.49496
R11739 iovss.n1160 iovss.n904 1.49496
R11740 iovss.n1149 iovss.n904 1.49496
R11741 iovss.n1217 iovss.n904 1.49494
R11742 iovss.n3090 iovss.n904 1.49489
R11743 iovss.n1172 iovss.n904 1.49489
R11744 iovss.n920 iovss.n904 1.49478
R11745 iovss.n1180 iovss.n904 1.49478
R11746 iovss.n1166 iovss.n904 1.49478
R11747 iovss.n1191 iovss.n904 1.49476
R11748 iovss.n1208 iovss.n904 1.49466
R11749 iovss.n3086 iovss.n904 1.49466
R11750 iovss.n1154 iovss.n904 1.49466
R11751 iovss.n1213 iovss.n904 1.49455
R11752 iovss.n918 iovss.n904 1.4945
R11753 iovss.n1209 iovss.n904 1.4945
R11754 iovss.n1146 iovss.n904 1.4945
R11755 iovss.n1174 iovss.n904 1.49432
R11756 iovss.n577 iovss.n571 1.10325
R11757 iovss.n2071 iovss.n2039 1.1005
R11758 iovss.n2070 iovss.n2040 1.1005
R11759 iovss.n2046 iovss.n2041 1.1005
R11760 iovss.n2061 iovss.n2047 1.1005
R11761 iovss.n2060 iovss.n2048 1.1005
R11762 iovss.n2059 iovss.n2049 1.1005
R11763 iovss.n2052 iovss.n2051 1.1005
R11764 iovss.n2050 iovss.n1508 1.1005
R11765 iovss.n2537 iovss.n1509 1.1005
R11766 iovss.n2536 iovss.n1510 1.1005
R11767 iovss.n2535 iovss.n1511 1.1005
R11768 iovss.n1517 iovss.n1512 1.1005
R11769 iovss.n2526 iovss.n1518 1.1005
R11770 iovss.n2525 iovss.n1519 1.1005
R11771 iovss.n2524 iovss.n1520 1.1005
R11772 iovss.n1525 iovss.n1521 1.1005
R11773 iovss.n2516 iovss.n1526 1.1005
R11774 iovss.n2515 iovss.n1527 1.1005
R11775 iovss.n2514 iovss.n1528 1.1005
R11776 iovss.n2406 iovss.n1529 1.1005
R11777 iovss.n2490 iovss.n2407 1.1005
R11778 iovss.n2489 iovss.n2408 1.1005
R11779 iovss.n2488 iovss.n2409 1.1005
R11780 iovss.n2430 iovss.n2410 1.1005
R11781 iovss.n2466 iovss.n2431 1.1005
R11782 iovss.n2465 iovss.n2432 1.1005
R11783 iovss.n2464 iovss.n2433 1.1005
R11784 iovss.n2435 iovss.n2434 1.1005
R11785 iovss.n1431 iovss.n1430 1.1005
R11786 iovss.n2591 iovss.n2590 1.1005
R11787 iovss.n2592 iovss.n1429 1.1005
R11788 iovss.n3463 iovss.n3462 1.1005
R11789 iovss.n3461 iovss.n63 1.1005
R11790 iovss.n3460 iovss.n3459 1.1005
R11791 iovss.n65 iovss.n64 1.1005
R11792 iovss.n3445 iovss.n73 1.1005
R11793 iovss.n3447 iovss.n3446 1.1005
R11794 iovss.n3444 iovss.n72 1.1005
R11795 iovss.n3443 iovss.n3442 1.1005
R11796 iovss.n75 iovss.n74 1.1005
R11797 iovss.n3318 iovss.n3317 1.1005
R11798 iovss.n3316 iovss.n464 1.1005
R11799 iovss.n3315 iovss.n3314 1.1005
R11800 iovss.n3312 iovss.n465 1.1005
R11801 iovss.n3310 iovss.n3308 1.1005
R11802 iovss.n3307 iovss.n467 1.1005
R11803 iovss.n3306 iovss.n3305 1.1005
R11804 iovss.n3303 iovss.n468 1.1005
R11805 iovss.n3301 iovss.n3299 1.1005
R11806 iovss.n3298 iovss.n469 1.1005
R11807 iovss.n3297 iovss.n3296 1.1005
R11808 iovss.n471 iovss.n470 1.1005
R11809 iovss.n3285 iovss.n3284 1.1005
R11810 iovss.n3283 iovss.n476 1.1005
R11811 iovss.n3282 iovss.n3281 1.1005
R11812 iovss.n478 iovss.n477 1.1005
R11813 iovss.n3269 iovss.n3268 1.1005
R11814 iovss.n3267 iovss.n483 1.1005
R11815 iovss.n3266 iovss.n3265 1.1005
R11816 iovss.n485 iovss.n484 1.1005
R11817 iovss.n604 iovss.n603 1.1005
R11818 iovss.n602 iovss.n563 1.1005
R11819 iovss.n601 iovss.n600 1.1005
R11820 iovss.n565 iovss.n564 1.1005
R11821 iovss.n590 iovss.n589 1.1005
R11822 iovss.n588 iovss.n570 1.1005
R11823 iovss.n587 iovss.n586 1.1005
R11824 iovss.n3464 iovss.n3463 1.1005
R11825 iovss.n63 iovss.n62 1.1005
R11826 iovss.n3459 iovss.n3458 1.1005
R11827 iovss.n3456 iovss.n65 1.1005
R11828 iovss.n73 iovss.n66 1.1005
R11829 iovss.n3448 iovss.n3447 1.1005
R11830 iovss.n72 iovss.n70 1.1005
R11831 iovss.n3442 iovss.n3441 1.1005
R11832 iovss.n76 iovss.n75 1.1005
R11833 iovss.n3319 iovss.n3318 1.1005
R11834 iovss.n464 iovss.n462 1.1005
R11835 iovss.n3314 iovss.n3313 1.1005
R11836 iovss.n3312 iovss.n3311 1.1005
R11837 iovss.n3310 iovss.n3309 1.1005
R11838 iovss.n467 iovss.n466 1.1005
R11839 iovss.n3305 iovss.n3304 1.1005
R11840 iovss.n3303 iovss.n3302 1.1005
R11841 iovss.n3301 iovss.n3300 1.1005
R11842 iovss.n3293 iovss.n469 1.1005
R11843 iovss.n3296 iovss.n3295 1.1005
R11844 iovss.n472 iovss.n471 1.1005
R11845 iovss.n3286 iovss.n3285 1.1005
R11846 iovss.n480 iovss.n476 1.1005
R11847 iovss.n3281 iovss.n3280 1.1005
R11848 iovss.n3271 iovss.n478 1.1005
R11849 iovss.n3270 iovss.n3269 1.1005
R11850 iovss.n487 iovss.n483 1.1005
R11851 iovss.n3265 iovss.n3264 1.1005
R11852 iovss.n561 iovss.n485 1.1005
R11853 iovss.n605 iovss.n604 1.1005
R11854 iovss.n563 iovss.n560 1.1005
R11855 iovss.n600 iovss.n599 1.1005
R11856 iovss.n566 iovss.n565 1.1005
R11857 iovss.n591 iovss.n590 1.1005
R11858 iovss.n574 iovss.n570 1.1005
R11859 iovss.n586 iovss.n585 1.1005
R11860 iovss.n575 iovss.n572 1.1005
R11861 iovss.n2177 iovss.n2161 0.826084
R11862 iovss.n776 iovss.n732 0.826084
R11863 iovss.n2342 iovss.n1223 0.822133
R11864 iovss.n3148 iovss.n884 0.822133
R11865 iovss.n3081 iovss.n1222 0.818682
R11866 iovss.n3082 iovss.n1221 0.818682
R11867 iovss.n1682 iovss.n1220 0.818682
R11868 iovss.n2351 iovss.n2350 0.818682
R11869 iovss.n2352 iovss.n1680 0.818682
R11870 iovss.n2353 iovss.n1679 0.818682
R11871 iovss.n2331 iovss.n1678 0.818682
R11872 iovss.n2329 iovss.n2328 0.818682
R11873 iovss.n2326 iovss.n2324 0.818682
R11874 iovss.n1689 iovss.n1688 0.818682
R11875 iovss.n2313 iovss.n2312 0.818682
R11876 iovss.n2310 iovss.n1693 0.818682
R11877 iovss.n2308 iovss.n2307 0.818682
R11878 iovss.n1697 iovss.n1696 0.818682
R11879 iovss.n2298 iovss.n2297 0.818682
R11880 iovss.n2295 iovss.n1701 0.818682
R11881 iovss.n2294 iovss.n1705 0.818682
R11882 iovss.n1881 iovss.n1703 0.818682
R11883 iovss.n2274 iovss.n2272 0.818682
R11884 iovss.n2276 iovss.n1879 0.818682
R11885 iovss.n2278 iovss.n1878 0.818682
R11886 iovss.n2280 iovss.n1877 0.818682
R11887 iovss.n2282 iovss.n1876 0.818682
R11888 iovss.n2284 iovss.n1875 0.818682
R11889 iovss.n2286 iovss.n1874 0.818682
R11890 iovss.n2287 iovss.n1873 0.818682
R11891 iovss.n2248 iovss.n1872 0.818682
R11892 iovss.n2246 iovss.n2245 0.818682
R11893 iovss.n2171 iovss.n1890 0.818682
R11894 iovss.n2202 iovss.n2200 0.818682
R11895 iovss.n2204 iovss.n2169 0.818682
R11896 iovss.n2178 iovss.n2163 0.818682
R11897 iovss.n2213 iovss.n2164 0.818682
R11898 iovss.n2212 iovss.n2165 0.818682
R11899 iovss.n2210 iovss.n2166 0.818682
R11900 iovss.n2208 iovss.n2167 0.818682
R11901 iovss.n2206 iovss.n2168 0.818682
R11902 iovss.n2935 iovss.n1223 0.818682
R11903 iovss.n3081 iovss.n3080 0.818682
R11904 iovss.n3083 iovss.n3082 0.818682
R11905 iovss.n1220 iovss.n1116 0.818682
R11906 iovss.n2351 iovss.n989 0.818682
R11907 iovss.n2352 iovss.n1677 0.818682
R11908 iovss.n2354 iovss.n2353 0.818682
R11909 iovss.n1678 iovss.n1653 0.818682
R11910 iovss.n2328 iovss.n2327 0.818682
R11911 iovss.n2326 iovss.n2325 0.818682
R11912 iovss.n1688 iovss.n1687 0.818682
R11913 iovss.n2312 iovss.n2311 0.818682
R11914 iovss.n2310 iovss.n2309 0.818682
R11915 iovss.n2308 iovss.n1593 0.818682
R11916 iovss.n1696 iovss.n1695 0.818682
R11917 iovss.n2297 iovss.n2296 0.818682
R11918 iovss.n2295 iovss.n1652 0.818682
R11919 iovss.n2294 iovss.n2293 0.818682
R11920 iovss.n1802 iovss.n1703 0.818682
R11921 iovss.n2274 iovss.n2273 0.818682
R11922 iovss.n2276 iovss.n2275 0.818682
R11923 iovss.n2278 iovss.n2277 0.818682
R11924 iovss.n2280 iovss.n2279 0.818682
R11925 iovss.n2282 iovss.n2281 0.818682
R11926 iovss.n2284 iovss.n2283 0.818682
R11927 iovss.n2286 iovss.n2285 0.818682
R11928 iovss.n2288 iovss.n2287 0.818682
R11929 iovss.n1872 iovss.n1871 0.818682
R11930 iovss.n2245 iovss.n2244 0.818682
R11931 iovss.n2100 iovss.n1890 0.818682
R11932 iovss.n2202 iovss.n2201 0.818682
R11933 iovss.n2204 iovss.n2203 0.818682
R11934 iovss.n2214 iovss.n2213 0.818682
R11935 iovss.n2212 iovss.n2211 0.818682
R11936 iovss.n2210 iovss.n2209 0.818682
R11937 iovss.n2208 iovss.n2207 0.818682
R11938 iovss.n2206 iovss.n2205 0.818682
R11939 iovss.n3164 iovss.n867 0.818682
R11940 iovss.n945 iovss.n868 0.818682
R11941 iovss.n3157 iovss.n875 0.818682
R11942 iovss.n3156 iovss.n876 0.818682
R11943 iovss.n914 iovss.n877 0.818682
R11944 iovss.n3149 iovss.n885 0.818682
R11945 iovss.n3148 iovss.n3147 0.818682
R11946 iovss.n3165 iovss.n866 0.818682
R11947 iovss.n859 iovss.n858 0.818682
R11948 iovss.n3172 iovss.n857 0.818682
R11949 iovss.n3173 iovss.n856 0.818682
R11950 iovss.n849 iovss.n848 0.818682
R11951 iovss.n3180 iovss.n847 0.818682
R11952 iovss.n3181 iovss.n245 0.818682
R11953 iovss.n840 iovss.n839 0.818682
R11954 iovss.n3188 iovss.n838 0.818682
R11955 iovss.n3189 iovss.n254 0.818682
R11956 iovss.n831 iovss.n276 0.818682
R11957 iovss.n3196 iovss.n830 0.818682
R11958 iovss.n3197 iovss.n829 0.818682
R11959 iovss.n822 iovss.n821 0.818682
R11960 iovss.n3204 iovss.n820 0.818682
R11961 iovss.n3205 iovss.n819 0.818682
R11962 iovss.n812 iovss.n811 0.818682
R11963 iovss.n3212 iovss.n810 0.818682
R11964 iovss.n3213 iovss.n809 0.818682
R11965 iovss.n802 iovss.n333 0.818682
R11966 iovss.n3220 iovss.n332 0.818682
R11967 iovss.n3221 iovss.n801 0.818682
R11968 iovss.n794 iovss.n793 0.818682
R11969 iovss.n3228 iovss.n792 0.818682
R11970 iovss.n3229 iovss.n791 0.818682
R11971 iovss.n784 iovss.n635 0.818682
R11972 iovss.n3236 iovss.n783 0.818682
R11973 iovss.n3237 iovss.n782 0.818682
R11974 iovss.n771 iovss.n770 0.818682
R11975 iovss.n3245 iovss.n3244 0.818682
R11976 iovss.n775 iovss.n769 0.818682
R11977 iovss.n3244 iovss.n3243 0.818682
R11978 iovss.n773 iovss.n771 0.818682
R11979 iovss.n3238 iovss.n3237 0.818682
R11980 iovss.n3236 iovss.n3235 0.818682
R11981 iovss.n785 iovss.n784 0.818682
R11982 iovss.n3230 iovss.n3229 0.818682
R11983 iovss.n3228 iovss.n3227 0.818682
R11984 iovss.n795 iovss.n794 0.818682
R11985 iovss.n3222 iovss.n3221 0.818682
R11986 iovss.n3220 iovss.n3219 0.818682
R11987 iovss.n803 iovss.n802 0.818682
R11988 iovss.n3214 iovss.n3213 0.818682
R11989 iovss.n3212 iovss.n3211 0.818682
R11990 iovss.n813 iovss.n812 0.818682
R11991 iovss.n3206 iovss.n3205 0.818682
R11992 iovss.n3204 iovss.n3203 0.818682
R11993 iovss.n823 iovss.n822 0.818682
R11994 iovss.n3198 iovss.n3197 0.818682
R11995 iovss.n3196 iovss.n3195 0.818682
R11996 iovss.n832 iovss.n831 0.818682
R11997 iovss.n3190 iovss.n3189 0.818682
R11998 iovss.n3188 iovss.n3187 0.818682
R11999 iovss.n841 iovss.n840 0.818682
R12000 iovss.n3182 iovss.n3181 0.818682
R12001 iovss.n3180 iovss.n3179 0.818682
R12002 iovss.n850 iovss.n849 0.818682
R12003 iovss.n3174 iovss.n3173 0.818682
R12004 iovss.n3172 iovss.n3171 0.818682
R12005 iovss.n860 iovss.n859 0.818682
R12006 iovss.n3166 iovss.n3165 0.818682
R12007 iovss.n3164 iovss.n3163 0.818682
R12008 iovss.n869 iovss.n868 0.818682
R12009 iovss.n3158 iovss.n3157 0.818682
R12010 iovss.n3156 iovss.n3155 0.818682
R12011 iovss.n878 iovss.n877 0.818682
R12012 iovss.n3150 iovss.n3149 0.818682
R12013 iovss.n2039 iovss.n2038 0.557177
R12014 iovss.n2593 iovss.n2592 0.557177
R12015 iovss.n587 iovss.n571 0.555375
R12016 iovss.n2897 iovss.n1249 0.541868
R12017 iovss.n2754 iovss.n2601 0.522214
R12018 iovss.n2765 iovss.n2763 0.452373
R12019 iovss.n2762 iovss.n2761 0.452373
R12020 iovss.n2241 iovss.n2161 0.414129
R12021 iovss.n3249 iovss.n732 0.414129
R12022 iovss.n1320 iovss 0.400946
R12023 iovss.n1319 iovss 0.400946
R12024 iovss.n3133 iovss 0.341436
R12025 iovss.n3362 iovss.n3344 0.302211
R12026 iovss.n3254 iovss.n3253 0.302211
R12027 iovss.n3432 iovss.n3431 0.302211
R12028 iovss.n46 iovss 0.301303
R12029 iovss.n3247 iovss.n3246 0.28175
R12030 iovss.n768 iovss.n767 0.28175
R12031 iovss.n756 iovss.n731 0.28175
R12032 iovss.n755 iovss.n657 0.28175
R12033 iovss.n754 iovss.n729 0.28175
R12034 iovss.n753 iovss.n658 0.28175
R12035 iovss.n752 iovss.n727 0.28175
R12036 iovss.n751 iovss.n659 0.28175
R12037 iovss.n750 iovss.n724 0.28175
R12038 iovss.n749 iovss.n660 0.28175
R12039 iovss.n748 iovss.n722 0.28175
R12040 iovss.n747 iovss.n661 0.28175
R12041 iovss.n746 iovss.n719 0.28175
R12042 iovss.n745 iovss.n662 0.28175
R12043 iovss.n744 iovss.n717 0.28175
R12044 iovss.n743 iovss.n663 0.28175
R12045 iovss.n714 iovss.n633 0.28175
R12046 iovss.n3252 iovss.n3251 0.28175
R12047 iovss.n712 iovss.n634 0.28175
R12048 iovss.n693 iovss.n664 0.28175
R12049 iovss.n710 iovss.n709 0.28175
R12050 iovss.n708 iovss.n665 0.28175
R12051 iovss.n707 iovss.n691 0.28175
R12052 iovss.n706 iovss.n666 0.28175
R12053 iovss.n705 iovss.n688 0.28175
R12054 iovss.n704 iovss.n667 0.28175
R12055 iovss.n703 iovss.n686 0.28175
R12056 iovss.n702 iovss.n668 0.28175
R12057 iovss.n701 iovss.n683 0.28175
R12058 iovss.n700 iovss.n669 0.28175
R12059 iovss.n699 iovss.n681 0.28175
R12060 iovss.n698 iovss.n670 0.28175
R12061 iovss.n697 iovss.n678 0.28175
R12062 iovss.n696 iovss.n671 0.28175
R12063 iovss.n695 iovss.n676 0.28175
R12064 iovss.n694 iovss.n672 0.28175
R12065 iovss.n3392 iovss.n334 0.28175
R12066 iovss.n359 iovss.n358 0.28175
R12067 iovss.n3390 iovss.n3389 0.28175
R12068 iovss.n3388 iovss.n3387 0.28175
R12069 iovss.n3377 iovss.n331 0.28175
R12070 iovss.n3376 iovss.n287 0.28175
R12071 iovss.n3375 iovss.n330 0.28175
R12072 iovss.n3374 iovss.n288 0.28175
R12073 iovss.n3373 iovss.n328 0.28175
R12074 iovss.n3372 iovss.n289 0.28175
R12075 iovss.n3371 iovss.n326 0.28175
R12076 iovss.n3370 iovss.n290 0.28175
R12077 iovss.n3369 iovss.n324 0.28175
R12078 iovss.n3368 iovss.n291 0.28175
R12079 iovss.n3367 iovss.n322 0.28175
R12080 iovss.n3366 iovss.n292 0.28175
R12081 iovss.n3365 iovss.n320 0.28175
R12082 iovss.n3364 iovss.n293 0.28175
R12083 iovss.n3363 iovss.n318 0.28175
R12084 iovss.n3361 iovss.n294 0.28175
R12085 iovss.n3360 iovss.n317 0.28175
R12086 iovss.n3359 iovss.n295 0.28175
R12087 iovss.n3358 iovss.n315 0.28175
R12088 iovss.n3357 iovss.n296 0.28175
R12089 iovss.n3356 iovss.n314 0.28175
R12090 iovss.n3355 iovss.n297 0.28175
R12091 iovss.n3354 iovss.n312 0.28175
R12092 iovss.n3353 iovss.n298 0.28175
R12093 iovss.n3352 iovss.n311 0.28175
R12094 iovss.n3351 iovss.n299 0.28175
R12095 iovss.n3350 iovss.n309 0.28175
R12096 iovss.n3349 iovss.n300 0.28175
R12097 iovss.n3348 iovss.n308 0.28175
R12098 iovss.n3347 iovss.n301 0.28175
R12099 iovss.n3346 iovss.n306 0.28175
R12100 iovss.n3345 iovss.n302 0.28175
R12101 iovss.n305 iovss.n264 0.28175
R12102 iovss.n3395 iovss.n3394 0.28175
R12103 iovss.n3427 iovss.n3413 0.28175
R12104 iovss.n3412 iovss.n263 0.28175
R12105 iovss.n3411 iovss.n253 0.28175
R12106 iovss.n3410 iovss.n203 0.28175
R12107 iovss.n3409 iovss.n251 0.28175
R12108 iovss.n3408 iovss.n204 0.28175
R12109 iovss.n3407 iovss.n250 0.28175
R12110 iovss.n3406 iovss.n205 0.28175
R12111 iovss.n3405 iovss.n248 0.28175
R12112 iovss.n3404 iovss.n206 0.28175
R12113 iovss.n3403 iovss.n247 0.28175
R12114 iovss.n3402 iovss.n207 0.28175
R12115 iovss.n3401 iovss.n245 0.28175
R12116 iovss.n3400 iovss.n208 0.28175
R12117 iovss.n3399 iovss.n243 0.28175
R12118 iovss.n3398 iovss.n209 0.28175
R12119 iovss.n3397 iovss.n241 0.28175
R12120 iovss.n3396 iovss.n210 0.28175
R12121 iovss.n239 iovss.n173 0.28175
R12122 iovss.n3430 iovss.n3429 0.28175
R12123 iovss.n237 iovss.n174 0.28175
R12124 iovss.n1321 iovss.n211 0.28175
R12125 iovss.n1322 iovss.n236 0.28175
R12126 iovss.n1323 iovss.n212 0.28175
R12127 iovss.n1324 iovss.n234 0.28175
R12128 iovss.n1325 iovss.n213 0.28175
R12129 iovss.n1326 iovss.n232 0.28175
R12130 iovss.n1327 iovss.n214 0.28175
R12131 iovss.n1328 iovss.n230 0.28175
R12132 iovss.n1329 iovss.n215 0.28175
R12133 iovss.n1330 iovss.n228 0.28175
R12134 iovss.n1331 iovss.n216 0.28175
R12135 iovss.n1332 iovss.n226 0.28175
R12136 iovss.n1333 iovss.n217 0.28175
R12137 iovss.n1334 iovss.n224 0.28175
R12138 iovss.n1335 iovss.n218 0.28175
R12139 iovss.n1336 iovss.n222 0.28175
R12140 iovss.n1337 iovss.n219 0.28175
R12141 iovss.n2177 iovss.n2176 0.201704
R12142 iovss.n777 iovss.n776 0.201704
R12143 iovss.n2343 iovss.n2342 0.2005
R12144 iovss.n2345 iovss.n2344 0.2005
R12145 iovss.n2347 iovss.n2346 0.2005
R12146 iovss.n2349 iovss.n2348 0.2005
R12147 iovss.n1683 iovss.n1681 0.2005
R12148 iovss.n2335 iovss.n2334 0.2005
R12149 iovss.n2333 iovss.n2332 0.2005
R12150 iovss.n2330 iovss.n1685 0.2005
R12151 iovss.n2321 iovss.n1686 0.2005
R12152 iovss.n2323 iovss.n2322 0.2005
R12153 iovss.n1694 iovss.n1690 0.2005
R12154 iovss.n2315 iovss.n2314 0.2005
R12155 iovss.n2306 iovss.n1692 0.2005
R12156 iovss.n2305 iovss.n2304 0.2005
R12157 iovss.n1702 iovss.n1698 0.2005
R12158 iovss.n2300 iovss.n2299 0.2005
R12159 iovss.n1704 iovss.n1700 0.2005
R12160 iovss.n2269 iovss.n2268 0.2005
R12161 iovss.n2271 iovss.n2270 0.2005
R12162 iovss.n1882 iovss.n1880 0.2005
R12163 iovss.n2263 iovss.n2262 0.2005
R12164 iovss.n2261 iovss.n2260 0.2005
R12165 iovss.n2259 iovss.n2258 0.2005
R12166 iovss.n1885 iovss.n1884 0.2005
R12167 iovss.n2254 iovss.n2253 0.2005
R12168 iovss.n2252 iovss.n2251 0.2005
R12169 iovss.n2250 iovss.n2249 0.2005
R12170 iovss.n2247 iovss.n1887 0.2005
R12171 iovss.n2197 iovss.n1889 0.2005
R12172 iovss.n2199 iovss.n2198 0.2005
R12173 iovss.n2172 iovss.n2170 0.2005
R12174 iovss.n2191 iovss.n2190 0.2005
R12175 iovss.n2189 iovss.n2188 0.2005
R12176 iovss.n2187 iovss.n2186 0.2005
R12177 iovss.n2175 iovss.n2174 0.2005
R12178 iovss.n2182 iovss.n2181 0.2005
R12179 iovss.n2180 iovss.n2179 0.2005
R12180 iovss.n884 iovss.n883 0.2005
R12181 iovss.n3152 iovss.n3151 0.2005
R12182 iovss.n3154 iovss.n3153 0.2005
R12183 iovss.n874 iovss.n873 0.2005
R12184 iovss.n3160 iovss.n3159 0.2005
R12185 iovss.n3162 iovss.n3161 0.2005
R12186 iovss.n865 iovss.n864 0.2005
R12187 iovss.n3168 iovss.n3167 0.2005
R12188 iovss.n3170 iovss.n3169 0.2005
R12189 iovss.n855 iovss.n854 0.2005
R12190 iovss.n3176 iovss.n3175 0.2005
R12191 iovss.n3178 iovss.n3177 0.2005
R12192 iovss.n846 iovss.n845 0.2005
R12193 iovss.n3184 iovss.n3183 0.2005
R12194 iovss.n3186 iovss.n3185 0.2005
R12195 iovss.n837 iovss.n836 0.2005
R12196 iovss.n3192 iovss.n3191 0.2005
R12197 iovss.n3194 iovss.n3193 0.2005
R12198 iovss.n828 iovss.n827 0.2005
R12199 iovss.n3200 iovss.n3199 0.2005
R12200 iovss.n3202 iovss.n3201 0.2005
R12201 iovss.n818 iovss.n817 0.2005
R12202 iovss.n3208 iovss.n3207 0.2005
R12203 iovss.n3210 iovss.n3209 0.2005
R12204 iovss.n808 iovss.n807 0.2005
R12205 iovss.n3216 iovss.n3215 0.2005
R12206 iovss.n3218 iovss.n3217 0.2005
R12207 iovss.n800 iovss.n799 0.2005
R12208 iovss.n3224 iovss.n3223 0.2005
R12209 iovss.n3226 iovss.n3225 0.2005
R12210 iovss.n790 iovss.n789 0.2005
R12211 iovss.n3232 iovss.n3231 0.2005
R12212 iovss.n3234 iovss.n3233 0.2005
R12213 iovss.n781 iovss.n780 0.2005
R12214 iovss.n3240 iovss.n3239 0.2005
R12215 iovss.n3242 iovss.n3241 0.2005
R12216 iovss.n774 iovss.n772 0.2005
R12217 iovss.n3248 iovss.n3247 0.144096
R12218 iovss.n3077 iovss 0.1105
R12219 iovss.n3107 iovss 0.1105
R12220 iovss.n1114 iovss 0.1105
R12221 iovss.n45 iovss 0.1105
R12222 iovss.n2343 iovss.n2341 0.1105
R12223 iovss.n2345 iovss.n2340 0.1105
R12224 iovss.n2347 iovss.n2339 0.1105
R12225 iovss.n2348 iovss.n2338 0.1105
R12226 iovss.n2337 iovss.n1683 0.1105
R12227 iovss.n2336 iovss.n2335 0.1105
R12228 iovss.n2333 iovss.n1684 0.1105
R12229 iovss.n2319 iovss.n1685 0.1105
R12230 iovss.n2321 iovss.n2320 0.1105
R12231 iovss.n2322 iovss.n2318 0.1105
R12232 iovss.n2317 iovss.n1690 0.1105
R12233 iovss.n2316 iovss.n2315 0.1105
R12234 iovss.n1692 iovss.n1691 0.1105
R12235 iovss.n2304 iovss.n2303 0.1105
R12236 iovss.n2302 iovss.n1698 0.1105
R12237 iovss.n2301 iovss.n2300 0.1105
R12238 iovss.n1700 iovss.n1699 0.1105
R12239 iovss.n2269 iovss.n2267 0.1105
R12240 iovss.n2270 iovss.n2266 0.1105
R12241 iovss.n2265 iovss.n1882 0.1105
R12242 iovss.n2264 iovss.n2263 0.1105
R12243 iovss.n2261 iovss.n1883 0.1105
R12244 iovss.n2259 iovss.n2257 0.1105
R12245 iovss.n2256 iovss.n1885 0.1105
R12246 iovss.n2255 iovss.n2254 0.1105
R12247 iovss.n2252 iovss.n1886 0.1105
R12248 iovss.n2250 iovss.n1888 0.1105
R12249 iovss.n2195 iovss.n1887 0.1105
R12250 iovss.n2197 iovss.n2196 0.1105
R12251 iovss.n2198 iovss.n2194 0.1105
R12252 iovss.n2193 iovss.n2172 0.1105
R12253 iovss.n2192 iovss.n2191 0.1105
R12254 iovss.n2189 iovss.n2173 0.1105
R12255 iovss.n2187 iovss.n2185 0.1105
R12256 iovss.n2184 iovss.n2175 0.1105
R12257 iovss.n2183 iovss.n2182 0.1105
R12258 iovss.n883 iovss.n882 0.1105
R12259 iovss.n3152 iovss.n881 0.1105
R12260 iovss.n3153 iovss.n880 0.1105
R12261 iovss.n879 iovss.n873 0.1105
R12262 iovss.n3160 iovss.n872 0.1105
R12263 iovss.n3161 iovss.n871 0.1105
R12264 iovss.n870 iovss.n864 0.1105
R12265 iovss.n3168 iovss.n863 0.1105
R12266 iovss.n3169 iovss.n862 0.1105
R12267 iovss.n861 iovss.n854 0.1105
R12268 iovss.n3176 iovss.n853 0.1105
R12269 iovss.n3177 iovss.n852 0.1105
R12270 iovss.n851 iovss.n845 0.1105
R12271 iovss.n3184 iovss.n844 0.1105
R12272 iovss.n3185 iovss.n843 0.1105
R12273 iovss.n842 iovss.n836 0.1105
R12274 iovss.n3192 iovss.n835 0.1105
R12275 iovss.n3193 iovss.n834 0.1105
R12276 iovss.n833 iovss.n827 0.1105
R12277 iovss.n3200 iovss.n826 0.1105
R12278 iovss.n3201 iovss.n825 0.1105
R12279 iovss.n824 iovss.n817 0.1105
R12280 iovss.n3208 iovss.n816 0.1105
R12281 iovss.n3209 iovss.n815 0.1105
R12282 iovss.n814 iovss.n807 0.1105
R12283 iovss.n3216 iovss.n806 0.1105
R12284 iovss.n3217 iovss.n805 0.1105
R12285 iovss.n804 iovss.n799 0.1105
R12286 iovss.n3224 iovss.n798 0.1105
R12287 iovss.n3225 iovss.n797 0.1105
R12288 iovss.n796 iovss.n789 0.1105
R12289 iovss.n3232 iovss.n788 0.1105
R12290 iovss.n3233 iovss.n787 0.1105
R12291 iovss.n786 iovss.n780 0.1105
R12292 iovss.n3240 iovss.n779 0.1105
R12293 iovss.n3241 iovss.n778 0.1105
R12294 iovss.n2073 iovss.n2034 0.0591667
R12295 iovss.n2073 iovss.n2037 0.0591667
R12296 iovss.n2069 iovss.n2037 0.0591667
R12297 iovss.n2069 iovss.n2042 0.0591667
R12298 iovss.n2062 iovss.n2042 0.0591667
R12299 iovss.n2062 iovss.n2045 0.0591667
R12300 iovss.n2058 iovss.n2045 0.0591667
R12301 iovss.n2058 iovss.n2053 0.0591667
R12302 iovss.n2053 iovss.n1506 0.0591667
R12303 iovss.n2538 iovss.n1506 0.0591667
R12304 iovss.n2538 iovss.n1507 0.0591667
R12305 iovss.n2534 iovss.n1507 0.0591667
R12306 iovss.n2534 iovss.n1513 0.0591667
R12307 iovss.n2527 iovss.n1513 0.0591667
R12308 iovss.n2527 iovss.n1516 0.0591667
R12309 iovss.n2523 iovss.n1516 0.0591667
R12310 iovss.n2523 iovss.n1522 0.0591667
R12311 iovss.n2517 iovss.n1522 0.0591667
R12312 iovss.n2517 iovss.n1524 0.0591667
R12313 iovss.n2513 iovss.n1524 0.0591667
R12314 iovss.n2513 iovss.n1530 0.0591667
R12315 iovss.n2491 iovss.n1530 0.0591667
R12316 iovss.n2491 iovss.n2405 0.0591667
R12317 iovss.n2487 iovss.n2405 0.0591667
R12318 iovss.n2487 iovss.n2411 0.0591667
R12319 iovss.n2467 iovss.n2411 0.0591667
R12320 iovss.n2467 iovss.n2429 0.0591667
R12321 iovss.n2463 iovss.n2429 0.0591667
R12322 iovss.n2463 iovss.n2436 0.0591667
R12323 iovss.n2436 iovss.n1432 0.0591667
R12324 iovss.n2589 iovss.n1432 0.0591667
R12325 iovss.n2589 iovss.n1427 0.0591667
R12326 iovss.n2595 iovss.n1427 0.0591667
R12327 iovss.n2595 iovss.n1428 0.0591667
R12328 iovss.n2076 iovss.n2075 0.0591667
R12329 iovss.n2075 iovss.n2036 0.0591667
R12330 iovss.n2068 iovss.n2036 0.0591667
R12331 iovss.n2068 iovss.n2066 0.0591667
R12332 iovss.n2066 iovss.n2064 0.0591667
R12333 iovss.n2064 iovss.n2044 0.0591667
R12334 iovss.n2057 iovss.n2044 0.0591667
R12335 iovss.n2057 iovss.n2055 0.0591667
R12336 iovss.n2055 iovss.n1503 0.0591667
R12337 iovss.n2539 iovss.n1503 0.0591667
R12338 iovss.n2539 iovss.n1505 0.0591667
R12339 iovss.n2533 iovss.n1505 0.0591667
R12340 iovss.n2533 iovss.n2531 0.0591667
R12341 iovss.n2531 iovss.n2529 0.0591667
R12342 iovss.n2529 iovss.n1515 0.0591667
R12343 iovss.n2522 iovss.n1515 0.0591667
R12344 iovss.n2522 iovss.n2520 0.0591667
R12345 iovss.n2520 iovss.n2519 0.0591667
R12346 iovss.n2519 iovss.n1523 0.0591667
R12347 iovss.n2512 iovss.n1523 0.0591667
R12348 iovss.n2512 iovss.n1531 0.0591667
R12349 iovss.n2492 iovss.n1531 0.0591667
R12350 iovss.n2492 iovss.n2404 0.0591667
R12351 iovss.n2486 iovss.n2404 0.0591667
R12352 iovss.n2486 iovss.n2412 0.0591667
R12353 iovss.n2468 iovss.n2412 0.0591667
R12354 iovss.n2468 iovss.n2428 0.0591667
R12355 iovss.n2462 iovss.n2428 0.0591667
R12356 iovss.n2462 iovss.n2437 0.0591667
R12357 iovss.n2437 iovss.n1433 0.0591667
R12358 iovss.n2588 iovss.n1433 0.0591667
R12359 iovss.n2588 iovss.n1414 0.0591667
R12360 iovss.n2596 iovss.n1414 0.0591667
R12361 iovss.n2596 iovss.n1426 0.0591667
R12362 iovss.n778 iovss.n777 0.0568704
R12363 iovss.n2183 iovss.n2176 0.0568704
R12364 iovss.n45 iovss 0.0555
R12365 iovss.n2965 iovss.n2964 0.0432778
R12366 iovss.n2966 iovss.n2965 0.0432778
R12367 iovss.n2967 iovss.n2966 0.0432778
R12368 iovss.n2968 iovss.n2967 0.0432778
R12369 iovss.n2969 iovss.n2968 0.0432778
R12370 iovss.n2970 iovss.n2969 0.0432778
R12371 iovss.n2971 iovss.n2970 0.0432778
R12372 iovss.n2972 iovss.n2971 0.0432778
R12373 iovss.n2973 iovss.n2972 0.0432778
R12374 iovss.n2974 iovss.n2973 0.0432778
R12375 iovss.n2974 iovss.n2960 0.0432778
R12376 iovss.n2980 iovss.n2960 0.0432778
R12377 iovss.n2981 iovss.n2980 0.0432778
R12378 iovss.n3068 iovss.n2981 0.0432778
R12379 iovss.n3068 iovss.n3067 0.0432778
R12380 iovss.n3067 iovss.n3065 0.0432778
R12381 iovss.n3065 iovss.n3063 0.0432778
R12382 iovss.n3063 iovss.n3061 0.0432778
R12383 iovss.n3061 iovss.n3059 0.0432778
R12384 iovss.n3059 iovss.n3057 0.0432778
R12385 iovss.n3057 iovss.n3055 0.0432778
R12386 iovss.n3055 iovss.n3053 0.0432778
R12387 iovss.n3053 iovss.n3051 0.0432778
R12388 iovss.n3051 iovss.n3049 0.0432778
R12389 iovss.n3049 iovss.n3047 0.0432778
R12390 iovss.n3047 iovss.n3045 0.0432778
R12391 iovss.n3045 iovss.n3043 0.0432778
R12392 iovss.n3043 iovss.n3041 0.0432778
R12393 iovss.n3041 iovss.n3039 0.0432778
R12394 iovss.n3039 iovss.n3037 0.0432778
R12395 iovss.n3037 iovss.n3035 0.0432778
R12396 iovss.n3035 iovss.n3033 0.0432778
R12397 iovss.n3033 iovss.n3031 0.0432778
R12398 iovss.n3031 iovss.n3029 0.0432778
R12399 iovss.n3029 iovss.n3027 0.0432778
R12400 iovss.n3027 iovss.n3025 0.0432778
R12401 iovss.n3025 iovss.n3023 0.0432778
R12402 iovss.n3023 iovss.n3021 0.0432778
R12403 iovss.n3021 iovss.n3019 0.0432778
R12404 iovss.n3019 iovss.n3017 0.0432778
R12405 iovss.n3017 iovss.n3015 0.0432778
R12406 iovss.n3015 iovss.n3013 0.0432778
R12407 iovss.n3013 iovss.n3011 0.0432778
R12408 iovss.n3011 iovss.n3009 0.0432778
R12409 iovss.n3009 iovss.n3007 0.0432778
R12410 iovss.n3007 iovss.n3005 0.0432778
R12411 iovss.n3005 iovss.n3003 0.0432778
R12412 iovss.n3003 iovss.n3001 0.0432778
R12413 iovss.n3001 iovss.n2999 0.0432778
R12414 iovss.n2999 iovss.n2997 0.0432778
R12415 iovss.n2997 iovss.n2995 0.0432778
R12416 iovss.n2995 iovss.n2993 0.0432778
R12417 iovss.n2993 iovss.n2991 0.0432778
R12418 iovss.n2991 iovss.n2989 0.0432778
R12419 iovss.n2989 iovss.n2987 0.0432778
R12420 iovss.n2987 iovss.n2985 0.0432778
R12421 iovss.n2985 iovss.n2983 0.0432778
R12422 iovss.n2983 iovss.n2933 0.0432778
R12423 iovss.n3073 iovss.n2933 0.0432778
R12424 iovss.n3074 iovss.n3073 0.0432778
R12425 iovss.n3075 iovss.n3074 0.0432778
R12426 iovss.n3128 iovss.n952 0.0432778
R12427 iovss.n3128 iovss.n3127 0.0432778
R12428 iovss.n3127 iovss.n3126 0.0432778
R12429 iovss.n3126 iovss.n3125 0.0432778
R12430 iovss.n3125 iovss.n3124 0.0432778
R12431 iovss.n3124 iovss.n3123 0.0432778
R12432 iovss.n3123 iovss.n3122 0.0432778
R12433 iovss.n3122 iovss.n3121 0.0432778
R12434 iovss.n3121 iovss.n3120 0.0432778
R12435 iovss.n3120 iovss.n953 0.0432778
R12436 iovss.n3116 iovss.n953 0.0432778
R12437 iovss.n3116 iovss.n3115 0.0432778
R12438 iovss.n3115 iovss.n3114 0.0432778
R12439 iovss.n3114 iovss.n958 0.0432778
R12440 iovss.n964 iovss.n958 0.0432778
R12441 iovss.n1058 iovss.n964 0.0432778
R12442 iovss.n1059 iovss.n1058 0.0432778
R12443 iovss.n1060 iovss.n1059 0.0432778
R12444 iovss.n1061 iovss.n1060 0.0432778
R12445 iovss.n1062 iovss.n1061 0.0432778
R12446 iovss.n1063 iovss.n1062 0.0432778
R12447 iovss.n1064 iovss.n1063 0.0432778
R12448 iovss.n1065 iovss.n1064 0.0432778
R12449 iovss.n1066 iovss.n1065 0.0432778
R12450 iovss.n1067 iovss.n1066 0.0432778
R12451 iovss.n1068 iovss.n1067 0.0432778
R12452 iovss.n1069 iovss.n1068 0.0432778
R12453 iovss.n1070 iovss.n1069 0.0432778
R12454 iovss.n1071 iovss.n1070 0.0432778
R12455 iovss.n1072 iovss.n1071 0.0432778
R12456 iovss.n1073 iovss.n1072 0.0432778
R12457 iovss.n1074 iovss.n1073 0.0432778
R12458 iovss.n1075 iovss.n1074 0.0432778
R12459 iovss.n1076 iovss.n1075 0.0432778
R12460 iovss.n1077 iovss.n1076 0.0432778
R12461 iovss.n1078 iovss.n1077 0.0432778
R12462 iovss.n1079 iovss.n1078 0.0432778
R12463 iovss.n1080 iovss.n1079 0.0432778
R12464 iovss.n1081 iovss.n1080 0.0432778
R12465 iovss.n1082 iovss.n1081 0.0432778
R12466 iovss.n1083 iovss.n1082 0.0432778
R12467 iovss.n1084 iovss.n1083 0.0432778
R12468 iovss.n1085 iovss.n1084 0.0432778
R12469 iovss.n1086 iovss.n1085 0.0432778
R12470 iovss.n1087 iovss.n1086 0.0432778
R12471 iovss.n1088 iovss.n1087 0.0432778
R12472 iovss.n1089 iovss.n1088 0.0432778
R12473 iovss.n1090 iovss.n1089 0.0432778
R12474 iovss.n1091 iovss.n1090 0.0432778
R12475 iovss.n1092 iovss.n1091 0.0432778
R12476 iovss.n1093 iovss.n1092 0.0432778
R12477 iovss.n1094 iovss.n1093 0.0432778
R12478 iovss.n1095 iovss.n1094 0.0432778
R12479 iovss.n1096 iovss.n1095 0.0432778
R12480 iovss.n1097 iovss.n1096 0.0432778
R12481 iovss.n1098 iovss.n1097 0.0432778
R12482 iovss.n1099 iovss.n1098 0.0432778
R12483 iovss.n1100 iovss.n1099 0.0432778
R12484 iovss.n1101 iovss.n1100 0.0432778
R12485 iovss.n1104 iovss.n1101 0.0432778
R12486 iovss.n1107 iovss.n1104 0.0432778
R12487 iovss.n2722 iovss.n2721 0.0347222
R12488 iovss.n2723 iovss.n2722 0.0347222
R12489 iovss.n2723 iovss.n2712 0.0347222
R12490 iovss.n2729 iovss.n2712 0.0347222
R12491 iovss.n2780 iovss.n2779 0.0347222
R12492 iovss.n2781 iovss.n2780 0.0347222
R12493 iovss.n2781 iovss.n1305 0.0347222
R12494 iovss.n2787 iovss.n1305 0.0347222
R12495 iovss.n2976 iovss.n2962 0.0347222
R12496 iovss.n2977 iovss.n2976 0.0347222
R12497 iovss.n2978 iovss.n2977 0.0347222
R12498 iovss.n2978 iovss.n2934 0.0347222
R12499 iovss.n1200 iovss.n1199 0.0347222
R12500 iovss.n1200 iovss.n1192 0.0347222
R12501 iovss.n1205 iovss.n1192 0.0347222
R12502 iovss.n1206 iovss.n1205 0.0347222
R12503 iovss.n955 iovss.n954 0.0347222
R12504 iovss.n956 iovss.n955 0.0347222
R12505 iovss.n959 iovss.n956 0.0347222
R12506 iovss.n960 iovss.n959 0.0347222
R12507 iovss.n3119 iovss.n938 0.0347222
R12508 iovss.n3119 iovss.n3118 0.0347222
R12509 iovss.n3118 iovss.n3117 0.0347222
R12510 iovss.n3117 iovss.n957 0.0347222
R12511 iovss.n3113 iovss.n957 0.0347222
R12512 iovss.n3113 iovss.n3112 0.0347222
R12513 iovss.n1106 iovss.n965 0.0347222
R12514 iovss.n1201 iovss.n1194 0.0347222
R12515 iovss.n1204 iovss.n1203 0.0347222
R12516 iovss.n3096 iovss.n1207 0.0347222
R12517 iovss.n2963 iovss.n892 0.0347222
R12518 iovss.n2975 iovss.n2963 0.0347222
R12519 iovss.n2975 iovss.n2961 0.0347222
R12520 iovss.n2979 iovss.n2961 0.0347222
R12521 iovss.n2979 iovss.n2959 0.0347222
R12522 iovss.n3069 iovss.n2959 0.0347222
R12523 iovss.n2778 iovss.n2776 0.0347222
R12524 iovss.n2778 iovss.n1307 0.0347222
R12525 iovss.n2782 iovss.n1307 0.0347222
R12526 iovss.n2784 iovss.n2782 0.0347222
R12527 iovss.n2786 iovss.n2784 0.0347222
R12528 iovss.n2786 iovss.n1225 0.0347222
R12529 iovss.n2720 iovss.n2718 0.0347222
R12530 iovss.n2720 iovss.n2714 0.0347222
R12531 iovss.n2724 iovss.n2714 0.0347222
R12532 iovss.n2726 iovss.n2724 0.0347222
R12533 iovss.n2728 iovss.n2726 0.0347222
R12534 iovss.n2728 iovss.n2711 0.0347222
R12535 iovss.n2762 iovss.n1337 0.0322121
R12536 iovss.n2685 iovss.n1365 0.0301825
R12537 iovss.n2828 iovss.n1263 0.0301825
R12538 iovss.n2619 iovss.n1364 0.0301477
R12539 iovss.n2826 iovss.n1262 0.0301477
R12540 iovss.n2757 iovss.n1351 0.0293095
R12541 iovss.n2609 iovss.n1390 0.0293095
R12542 iovss.n2627 iovss.n1398 0.0293095
R12543 iovss.n2643 iovss.n1352 0.0293095
R12544 iovss.n1315 iovss.n1276 0.0293095
R12545 iovss.n2801 iovss.n1288 0.0293095
R12546 iovss.n2846 iovss.n1296 0.0293095
R12547 iovss.n2890 iovss.n1250 0.0293095
R12548 iovss.n2725 iovss.n1374 0.0284365
R12549 iovss.n2709 iovss.n1386 0.0284365
R12550 iovss.n2661 iovss.n1402 0.0284365
R12551 iovss.n2658 iovss.n1356 0.0284365
R12552 iovss.n2783 iovss.n1272 0.0284365
R12553 iovss.n1284 iovss.n1283 0.0284365
R12554 iovss.n2868 iovss.n1300 0.0284365
R12555 iovss.n2873 iovss.n1254 0.0284365
R12556 iovss.n1320 iovss.t5 0.0282811
R12557 iovss.n1319 iovss.t4 0.0282811
R12558 iovss.n1378 iovss.n1377 0.0280247
R12559 iovss.n2700 iovss.n1370 0.0280247
R12560 iovss.n2670 iovss.n1399 0.0280247
R12561 iovss.n2649 iovss.n1406 0.0280247
R12562 iovss.n2770 iovss.n1275 0.0280247
R12563 iovss.n2803 iovss.n1268 0.0280247
R12564 iovss.n2853 iovss.n1297 0.0280247
R12565 iovss.n2891 iovss.n1304 0.0280247
R12566 iovss.n1350 iovss.n1349 0.0275635
R12567 iovss.n2611 iovss.n1369 0.0275635
R12568 iovss.n2625 iovss.n1361 0.0275635
R12569 iovss.n1408 iovss.n1407 0.0275635
R12570 iovss.n1317 iovss.n1278 0.0275635
R12571 iovss.n2806 iovss.n1267 0.0275635
R12572 iovss.n2841 iovss.n1259 0.0275635
R12573 iovss.n2894 iovss.n1248 0.0275635
R12574 iovss.n2715 iovss.n1385 0.0271517
R12575 iovss.n2603 iovss.n1387 0.0271517
R12576 iovss.n2633 iovss.n1357 0.0271517
R12577 iovss.n2637 iovss.n1355 0.0271517
R12578 iovss.n1308 iovss.n1282 0.0271517
R12579 iovss.n2788 iovss.n1285 0.0271517
R12580 iovss.n2861 iovss.n1255 0.0271517
R12581 iovss.n2871 iovss.n1253 0.0271517
R12582 iovss.n2688 iovss.n1393 0.0266905
R12583 iovss.n2682 iovss.n1394 0.0266905
R12584 iovss.n2823 iovss.n1291 0.0266905
R12585 iovss.n2833 iovss.n1292 0.0266905
R12586 iovss.n2694 iovss.n1368 0.0262787
R12587 iovss.n2676 iovss.n1397 0.0262787
R12588 iovss.n2756 iovss.n2755 0.0262787
R12589 iovss.n2813 iovss.n1266 0.0262787
R12590 iovss.n2843 iovss.n1295 0.0262787
R12591 iovss.n2896 iovss.n2895 0.0262787
R12592 iovss.n1382 iovss.n1379 0.0258175
R12593 iovss.n2607 iovss.n1371 0.0258175
R12594 iovss.n2629 iovss.n1360 0.0258175
R12595 iovss.n2641 iovss.n1405 0.0258175
R12596 iovss.n1314 iovss.n1279 0.0258175
R12597 iovss.n2796 iovss.n1269 0.0258175
R12598 iovss.n2851 iovss.n1258 0.0258175
R12599 iovss.n2881 iovss.n1303 0.0258175
R12600 iovss.n2615 iovss.n1366 0.0254057
R12601 iovss.n2621 iovss.n1395 0.0254057
R12602 iovss.n2816 iovss.n1264 0.0254057
R12603 iovss.n2831 iovss.n1293 0.0254057
R12604 iovss.n2713 iovss.n1384 0.0249444
R12605 iovss.n2706 iovss.n1373 0.0249444
R12606 iovss.n2664 iovss.n1358 0.0249444
R12607 iovss.n2655 iovss.n1403 0.0249444
R12608 iovss.n1306 iovss.n1281 0.0249444
R12609 iovss.n2793 iovss.n1271 0.0249444
R12610 iovss.n2863 iovss.n1256 0.0249444
R12611 iovss.n2878 iovss.n1301 0.0249444
R12612 iovss.n2717 iovss.n1383 0.0245327
R12613 iovss.n2703 iovss.n1389 0.0245327
R12614 iovss.n2667 iovss.n1359 0.0245327
R12615 iovss.n2652 iovss.n1353 0.0245327
R12616 iovss.n1311 iovss.n1280 0.0245327
R12617 iovss.n2798 iovss.n1287 0.0245327
R12618 iovss.n2858 iovss.n1257 0.0245327
R12619 iovss.n2883 iovss.n1251 0.0245327
R12620 iovss.n2613 iovss.n1391 0.0240714
R12621 iovss.n2623 iovss.n1396 0.0240714
R12622 iovss.n2811 iovss.n1289 0.0240714
R12623 iovss.n2836 iovss.n1294 0.0240714
R12624 iovss.n2719 iovss.n1375 0.0236596
R12625 iovss.n2605 iovss.n1372 0.0236596
R12626 iovss.n2631 iovss.n1401 0.0236596
R12627 iovss.n2639 iovss.n1404 0.0236596
R12628 iovss.n2777 iovss.n1273 0.0236596
R12629 iovss.n2791 iovss.n1270 0.0236596
R12630 iovss.n2856 iovss.n1299 0.0236596
R12631 iovss.n2876 iovss.n1302 0.0236596
R12632 iovss.n2691 iovss.n1367 0.0231984
R12633 iovss.n2679 iovss.n1363 0.0231984
R12634 iovss.n2818 iovss.n1265 0.0231984
R12635 iovss.n2838 iovss.n1261 0.0231984
R12636 iovss.n2964 iovss.n904 0.0231984
R12637 iovss.n952 iovss.n904 0.0231984
R12638 iovss.n2691 iovss.n1392 0.0227866
R12639 iovss.n2679 iovss.n1362 0.0227866
R12640 iovss.n2818 iovss.n1290 0.0227866
R12641 iovss.n2838 iovss.n1260 0.0227866
R12642 iovss.n581 iovss.n579 0.0225
R12643 iovss.n583 iovss.n581 0.0225
R12644 iovss.n583 iovss.n568 0.0225
R12645 iovss.n594 iovss.n568 0.0225
R12646 iovss.n596 iovss.n594 0.0225
R12647 iovss.n596 iovss.n559 0.0225
R12648 iovss.n607 iovss.n559 0.0225
R12649 iovss.n607 iovss.n488 0.0225
R12650 iovss.n3261 iovss.n488 0.0225
R12651 iovss.n3262 iovss.n3261 0.0225
R12652 iovss.n3262 iovss.n481 0.0225
R12653 iovss.n3274 iovss.n481 0.0225
R12654 iovss.n3276 iovss.n3274 0.0225
R12655 iovss.n3278 iovss.n3276 0.0225
R12656 iovss.n3278 iovss.n474 0.0225
R12657 iovss.n3289 iovss.n474 0.0225
R12658 iovss.n3291 iovss.n3289 0.0225
R12659 iovss.n3291 iovss.n453 0.0225
R12660 iovss.n3337 iovss.n453 0.0225
R12661 iovss.n3337 iovss.n3336 0.0225
R12662 iovss.n3336 iovss.n3332 0.0225
R12663 iovss.n3332 iovss.n3331 0.0225
R12664 iovss.n3331 iovss.n3329 0.0225
R12665 iovss.n3329 iovss.n3327 0.0225
R12666 iovss.n3327 iovss.n3326 0.0225
R12667 iovss.n3326 iovss.n3324 0.0225
R12668 iovss.n3324 iovss.n3322 0.0225
R12669 iovss.n3322 iovss.n77 0.0225
R12670 iovss.n3438 iovss.n77 0.0225
R12671 iovss.n3438 iovss.n69 0.0225
R12672 iovss.n3450 iovss.n69 0.0225
R12673 iovss.n3450 iovss.n67 0.0225
R12674 iovss.n3454 iovss.n67 0.0225
R12675 iovss.n3454 iovss.n59 0.0225
R12676 iovss.n3469 iovss.n59 0.0225
R12677 iovss.n3469 iovss.n3468 0.0225
R12678 iovss.n3468 iovss.n3466 0.0225
R12679 iovss.n3335 iovss.n3334 0.0225
R12680 iovss.n3452 iovss.n3451 0.0225
R12681 iovss.n3453 iovss.n3452 0.0225
R12682 iovss.n3453 iovss.n58 0.0225
R12683 iovss.n3470 iovss.n58 0.0225
R12684 iovss.n2719 iovss.n1376 0.0223254
R12685 iovss.n2605 iovss.n1388 0.0223254
R12686 iovss.n2631 iovss.n1400 0.0223254
R12687 iovss.n2639 iovss.n1354 0.0223254
R12688 iovss.n2777 iovss.n1274 0.0223254
R12689 iovss.n2791 iovss.n1286 0.0223254
R12690 iovss.n2856 iovss.n1298 0.0223254
R12691 iovss.n2876 iovss.n1252 0.0223254
R12692 iovss.n2242 iovss.n2093 0.0220831
R12693 iovss.n2291 iovss.n1502 0.0220831
R12694 iovss.n2398 iovss.n2397 0.0220831
R12695 iovss.n2613 iovss.n1392 0.0219136
R12696 iovss.n2623 iovss.n1362 0.0219136
R12697 iovss.n2811 iovss.n1290 0.0219136
R12698 iovss.n2836 iovss.n1260 0.0219136
R12699 iovss.n2763 iovss.n2762 0.0217675
R12700 iovss.n2717 iovss.n1376 0.0214524
R12701 iovss.n2703 iovss.n1388 0.0214524
R12702 iovss.n2667 iovss.n1400 0.0214524
R12703 iovss.n2652 iovss.n1354 0.0214524
R12704 iovss.n1311 iovss.n1274 0.0214524
R12705 iovss.n2798 iovss.n1286 0.0214524
R12706 iovss.n2858 iovss.n1298 0.0214524
R12707 iovss.n2883 iovss.n1252 0.0214524
R12708 iovss.n2713 iovss.n1375 0.0210406
R12709 iovss.n2706 iovss.n1372 0.0210406
R12710 iovss.n2664 iovss.n1401 0.0210406
R12711 iovss.n2655 iovss.n1404 0.0210406
R12712 iovss.n1306 iovss.n1273 0.0210406
R12713 iovss.n2793 iovss.n1270 0.0210406
R12714 iovss.n2863 iovss.n1299 0.0210406
R12715 iovss.n2878 iovss.n1302 0.0210406
R12716 iovss.n2615 iovss.n1367 0.0205794
R12717 iovss.n2621 iovss.n1363 0.0205794
R12718 iovss.n2816 iovss.n1265 0.0205794
R12719 iovss.n2831 iovss.n1261 0.0205794
R12720 iovss.n927 iovss.n904 0.0205794
R12721 iovss.n3132 iovss.n904 0.0205794
R12722 iovss.n1383 iovss.n1382 0.0201676
R12723 iovss.n2607 iovss.n1389 0.0201676
R12724 iovss.n2629 iovss.n1359 0.0201676
R12725 iovss.n2641 iovss.n1353 0.0201676
R12726 iovss.n1314 iovss.n1280 0.0201676
R12727 iovss.n2796 iovss.n1287 0.0201676
R12728 iovss.n2851 iovss.n1257 0.0201676
R12729 iovss.n2881 iovss.n1251 0.0201676
R12730 iovss.n3451 iovss.n68 0.01975
R12731 iovss.n2694 iovss.n1391 0.0197063
R12732 iovss.n2676 iovss.n1396 0.0197063
R12733 iovss.n2813 iovss.n1289 0.0197063
R12734 iovss.n2843 iovss.n1294 0.0197063
R12735 iovss.n2688 iovss.n1366 0.0192946
R12736 iovss.n2682 iovss.n1395 0.0192946
R12737 iovss.n2823 iovss.n1264 0.0192946
R12738 iovss.n2833 iovss.n1293 0.0192946
R12739 iovss.n2715 iovss.n1384 0.0188333
R12740 iovss.n2603 iovss.n1373 0.0188333
R12741 iovss.n2633 iovss.n1358 0.0188333
R12742 iovss.n2637 iovss.n1403 0.0188333
R12743 iovss.n1308 iovss.n1281 0.0188333
R12744 iovss.n2788 iovss.n1271 0.0188333
R12745 iovss.n2861 iovss.n1256 0.0188333
R12746 iovss.n2871 iovss.n1301 0.0188333
R12747 iovss.n1349 iovss.n1339 0.0187533
R12748 iovss.n1317 iovss.n1277 0.0187533
R12749 iovss.n3343 iovss.n380 0.01865
R12750 iovss.n2611 iovss.n1368 0.0184215
R12751 iovss.n2625 iovss.n1397 0.0184215
R12752 iovss.n2756 iovss.n1408 0.0184215
R12753 iovss.n2806 iovss.n1266 0.0184215
R12754 iovss.n2841 iovss.n1295 0.0184215
R12755 iovss.n2895 iovss.n1248 0.0184215
R12756 iovss.n933 iovss.n931 0.0180786
R12757 iovss.n3131 iovss.n928 0.0180786
R12758 iovss.n934 iovss.n929 0.0180786
R12759 iovss.n3129 iovss.n950 0.0180786
R12760 iovss.n951 iovss.n935 0.0180786
R12761 iovss.n948 iovss.n944 0.0180786
R12762 iovss.n943 iovss.n936 0.0180786
R12763 iovss.n947 iovss.n942 0.0180786
R12764 iovss.n941 iovss.n937 0.0180786
R12765 iovss.n946 iovss.n940 0.0180786
R12766 iovss.n939 iovss.n938 0.0180786
R12767 iovss.n3111 iovss.n3110 0.0180786
R12768 iovss.n1033 iovss.n963 0.0180786
R12769 iovss.n1032 iovss.n966 0.0180786
R12770 iovss.n1055 iovss.n1031 0.0180786
R12771 iovss.n1030 iovss.n967 0.0180786
R12772 iovss.n1054 iovss.n1029 0.0180786
R12773 iovss.n1028 iovss.n968 0.0180786
R12774 iovss.n1053 iovss.n1027 0.0180786
R12775 iovss.n1026 iovss.n969 0.0180786
R12776 iovss.n1052 iovss.n1025 0.0180786
R12777 iovss.n1024 iovss.n970 0.0180786
R12778 iovss.n1051 iovss.n1023 0.0180786
R12779 iovss.n1022 iovss.n971 0.0180786
R12780 iovss.n1050 iovss.n1021 0.0180786
R12781 iovss.n1020 iovss.n972 0.0180786
R12782 iovss.n1049 iovss.n1019 0.0180786
R12783 iovss.n1018 iovss.n973 0.0180786
R12784 iovss.n1048 iovss.n1017 0.0180786
R12785 iovss.n1016 iovss.n974 0.0180786
R12786 iovss.n1047 iovss.n1015 0.0180786
R12787 iovss.n1014 iovss.n975 0.0180786
R12788 iovss.n1046 iovss.n1013 0.0180786
R12789 iovss.n1012 iovss.n976 0.0180786
R12790 iovss.n1045 iovss.n1011 0.0180786
R12791 iovss.n1010 iovss.n977 0.0180786
R12792 iovss.n1044 iovss.n1009 0.0180786
R12793 iovss.n1008 iovss.n978 0.0180786
R12794 iovss.n1043 iovss.n1007 0.0180786
R12795 iovss.n1006 iovss.n979 0.0180786
R12796 iovss.n1042 iovss.n1005 0.0180786
R12797 iovss.n1004 iovss.n980 0.0180786
R12798 iovss.n1041 iovss.n1003 0.0180786
R12799 iovss.n1002 iovss.n981 0.0180786
R12800 iovss.n1040 iovss.n1001 0.0180786
R12801 iovss.n1000 iovss.n982 0.0180786
R12802 iovss.n1039 iovss.n999 0.0180786
R12803 iovss.n998 iovss.n983 0.0180786
R12804 iovss.n1038 iovss.n997 0.0180786
R12805 iovss.n996 iovss.n984 0.0180786
R12806 iovss.n1037 iovss.n995 0.0180786
R12807 iovss.n994 iovss.n985 0.0180786
R12808 iovss.n1036 iovss.n993 0.0180786
R12809 iovss.n992 iovss.n986 0.0180786
R12810 iovss.n1035 iovss.n991 0.0180786
R12811 iovss.n990 iovss.n987 0.0180786
R12812 iovss.n1103 iovss.n1102 0.0180786
R12813 iovss.n1106 iovss.n988 0.0180786
R12814 iovss.n3108 iovss.n1034 0.0180786
R12815 iovss.n908 iovss.n906 0.0180786
R12816 iovss.n3135 iovss.n925 0.0180786
R12817 iovss.n926 iovss.n909 0.0180786
R12818 iovss.n1195 iovss.n910 0.0180786
R12819 iovss.n921 iovss.n911 0.0180786
R12820 iovss.n1197 iovss.n919 0.0180786
R12821 iovss.n916 iovss.n915 0.0180786
R12822 iovss.n1196 iovss.n913 0.0180786
R12823 iovss.n1190 iovss.n1188 0.0180786
R12824 iovss.n1187 iovss.n1185 0.0180786
R12825 iovss.n1184 iovss.n1183 0.0180786
R12826 iovss.n3093 iovss.n1182 0.0180786
R12827 iovss.n3092 iovss.n1120 0.0180786
R12828 iovss.n1179 iovss.n1121 0.0180786
R12829 iovss.n1177 iovss.n1122 0.0180786
R12830 iovss.n1212 iovss.n1123 0.0180786
R12831 iovss.n1211 iovss.n1175 0.0180786
R12832 iovss.n1173 iovss.n1171 0.0180786
R12833 iovss.n1170 iovss.n1168 0.0180786
R12834 iovss.n1167 iovss.n1165 0.0180786
R12835 iovss.n1164 iovss.n1163 0.0180786
R12836 iovss.n3089 iovss.n1162 0.0180786
R12837 iovss.n3088 iovss.n1128 0.0180786
R12838 iovss.n1159 iovss.n1129 0.0180786
R12839 iovss.n1157 iovss.n1130 0.0180786
R12840 iovss.n1216 iovss.n1131 0.0180786
R12841 iovss.n1215 iovss.n1155 0.0180786
R12842 iovss.n1153 iovss.n1151 0.0180786
R12843 iovss.n1150 iovss.n1148 0.0180786
R12844 iovss.n1147 iovss.n1145 0.0180786
R12845 iovss.n1144 iovss.n1143 0.0180786
R12846 iovss.n3085 iovss.n1142 0.0180786
R12847 iovss.n3084 iovss.n1136 0.0180786
R12848 iovss.n1139 iovss.n1138 0.0180786
R12849 iovss.n1138 iovss.n1109 0.0180786
R12850 iovss.n3099 iovss.n1108 0.0180786
R12851 iovss.n1034 iovss.n965 0.0180786
R12852 iovss.n903 iovss.n887 0.0180786
R12853 iovss.n3143 iovss.n902 0.0180786
R12854 iovss.n901 iovss.n888 0.0180786
R12855 iovss.n3142 iovss.n900 0.0180786
R12856 iovss.n899 iovss.n889 0.0180786
R12857 iovss.n3141 iovss.n898 0.0180786
R12858 iovss.n897 iovss.n890 0.0180786
R12859 iovss.n3140 iovss.n896 0.0180786
R12860 iovss.n895 iovss.n891 0.0180786
R12861 iovss.n3139 iovss.n894 0.0180786
R12862 iovss.n893 iovss.n892 0.0180786
R12863 iovss.n3066 iovss.n2902 0.0180786
R12864 iovss.n3064 iovss.n2958 0.0180786
R12865 iovss.n3062 iovss.n2903 0.0180786
R12866 iovss.n3060 iovss.n2957 0.0180786
R12867 iovss.n3058 iovss.n2904 0.0180786
R12868 iovss.n3056 iovss.n2956 0.0180786
R12869 iovss.n3054 iovss.n2905 0.0180786
R12870 iovss.n3052 iovss.n2955 0.0180786
R12871 iovss.n3050 iovss.n2906 0.0180786
R12872 iovss.n3048 iovss.n2954 0.0180786
R12873 iovss.n3046 iovss.n2907 0.0180786
R12874 iovss.n3044 iovss.n2953 0.0180786
R12875 iovss.n3042 iovss.n2908 0.0180786
R12876 iovss.n3040 iovss.n2952 0.0180786
R12877 iovss.n3038 iovss.n2909 0.0180786
R12878 iovss.n3036 iovss.n2951 0.0180786
R12879 iovss.n3034 iovss.n2910 0.0180786
R12880 iovss.n3032 iovss.n2950 0.0180786
R12881 iovss.n3030 iovss.n2911 0.0180786
R12882 iovss.n3028 iovss.n2949 0.0180786
R12883 iovss.n3026 iovss.n2912 0.0180786
R12884 iovss.n3024 iovss.n2948 0.0180786
R12885 iovss.n3022 iovss.n2913 0.0180786
R12886 iovss.n3020 iovss.n2947 0.0180786
R12887 iovss.n3018 iovss.n2914 0.0180786
R12888 iovss.n3016 iovss.n2946 0.0180786
R12889 iovss.n3014 iovss.n2915 0.0180786
R12890 iovss.n3012 iovss.n2945 0.0180786
R12891 iovss.n3010 iovss.n2916 0.0180786
R12892 iovss.n3008 iovss.n2944 0.0180786
R12893 iovss.n3006 iovss.n2917 0.0180786
R12894 iovss.n3004 iovss.n2943 0.0180786
R12895 iovss.n3002 iovss.n2918 0.0180786
R12896 iovss.n3000 iovss.n2942 0.0180786
R12897 iovss.n2998 iovss.n2919 0.0180786
R12898 iovss.n2996 iovss.n2941 0.0180786
R12899 iovss.n2994 iovss.n2920 0.0180786
R12900 iovss.n2992 iovss.n2940 0.0180786
R12901 iovss.n2990 iovss.n2921 0.0180786
R12902 iovss.n2988 iovss.n2939 0.0180786
R12903 iovss.n2986 iovss.n2922 0.0180786
R12904 iovss.n2984 iovss.n2938 0.0180786
R12905 iovss.n2982 iovss.n2923 0.0180786
R12906 iovss.n2937 iovss.n2936 0.0180786
R12907 iovss.n3072 iovss.n2924 0.0180786
R12908 iovss.n3071 iovss.n2926 0.0180786
R12909 iovss.n2928 iovss.n2925 0.0180786
R12910 iovss.n3078 iovss.n2927 0.0180786
R12911 iovss.n3078 iovss.n2932 0.0180786
R12912 iovss.n3076 iovss.n2932 0.0180786
R12913 iovss.n2927 iovss.n2925 0.0180786
R12914 iovss.n2928 iovss.n2926 0.0180786
R12915 iovss.n3072 iovss.n3071 0.0180786
R12916 iovss.n2936 iovss.n2924 0.0180786
R12917 iovss.n2982 iovss.n2937 0.0180786
R12918 iovss.n2984 iovss.n2923 0.0180786
R12919 iovss.n2986 iovss.n2938 0.0180786
R12920 iovss.n2988 iovss.n2922 0.0180786
R12921 iovss.n2990 iovss.n2939 0.0180786
R12922 iovss.n2992 iovss.n2921 0.0180786
R12923 iovss.n2994 iovss.n2940 0.0180786
R12924 iovss.n2996 iovss.n2920 0.0180786
R12925 iovss.n2998 iovss.n2941 0.0180786
R12926 iovss.n3000 iovss.n2919 0.0180786
R12927 iovss.n3002 iovss.n2942 0.0180786
R12928 iovss.n3004 iovss.n2918 0.0180786
R12929 iovss.n3006 iovss.n2943 0.0180786
R12930 iovss.n3008 iovss.n2917 0.0180786
R12931 iovss.n3010 iovss.n2944 0.0180786
R12932 iovss.n3012 iovss.n2916 0.0180786
R12933 iovss.n3014 iovss.n2945 0.0180786
R12934 iovss.n3016 iovss.n2915 0.0180786
R12935 iovss.n3018 iovss.n2946 0.0180786
R12936 iovss.n3020 iovss.n2914 0.0180786
R12937 iovss.n3022 iovss.n2947 0.0180786
R12938 iovss.n3024 iovss.n2913 0.0180786
R12939 iovss.n3026 iovss.n2948 0.0180786
R12940 iovss.n3028 iovss.n2912 0.0180786
R12941 iovss.n3030 iovss.n2949 0.0180786
R12942 iovss.n3032 iovss.n2911 0.0180786
R12943 iovss.n3034 iovss.n2950 0.0180786
R12944 iovss.n3036 iovss.n2910 0.0180786
R12945 iovss.n3038 iovss.n2951 0.0180786
R12946 iovss.n3040 iovss.n2909 0.0180786
R12947 iovss.n3042 iovss.n2952 0.0180786
R12948 iovss.n3044 iovss.n2908 0.0180786
R12949 iovss.n3046 iovss.n2953 0.0180786
R12950 iovss.n3048 iovss.n2907 0.0180786
R12951 iovss.n3050 iovss.n2954 0.0180786
R12952 iovss.n3052 iovss.n2906 0.0180786
R12953 iovss.n3054 iovss.n2955 0.0180786
R12954 iovss.n3056 iovss.n2905 0.0180786
R12955 iovss.n3058 iovss.n2956 0.0180786
R12956 iovss.n3060 iovss.n2904 0.0180786
R12957 iovss.n3062 iovss.n2957 0.0180786
R12958 iovss.n3064 iovss.n2903 0.0180786
R12959 iovss.n3066 iovss.n2958 0.0180786
R12960 iovss.n3069 iovss.n2902 0.0180786
R12961 iovss.n1141 iovss.n1139 0.0180786
R12962 iovss.n3085 iovss.n3084 0.0180786
R12963 iovss.n1218 iovss.n1142 0.0180786
R12964 iovss.n1143 iovss.n1135 0.0180786
R12965 iovss.n1145 iovss.n1134 0.0180786
R12966 iovss.n1148 iovss.n1133 0.0180786
R12967 iovss.n1151 iovss.n1132 0.0180786
R12968 iovss.n1216 iovss.n1215 0.0180786
R12969 iovss.n3087 iovss.n1131 0.0180786
R12970 iovss.n1158 iovss.n1157 0.0180786
R12971 iovss.n1161 iovss.n1159 0.0180786
R12972 iovss.n3089 iovss.n3088 0.0180786
R12973 iovss.n1214 iovss.n1162 0.0180786
R12974 iovss.n1163 iovss.n1127 0.0180786
R12975 iovss.n1165 iovss.n1126 0.0180786
R12976 iovss.n1168 iovss.n1125 0.0180786
R12977 iovss.n1171 iovss.n1124 0.0180786
R12978 iovss.n1212 iovss.n1211 0.0180786
R12979 iovss.n3091 iovss.n1123 0.0180786
R12980 iovss.n1178 iovss.n1177 0.0180786
R12981 iovss.n1181 iovss.n1179 0.0180786
R12982 iovss.n3093 iovss.n3092 0.0180786
R12983 iovss.n1210 iovss.n1182 0.0180786
R12984 iovss.n1183 iovss.n1119 0.0180786
R12985 iovss.n1185 iovss.n1118 0.0180786
R12986 iovss.n1188 iovss.n1117 0.0180786
R12987 iovss.n3100 iovss.n1109 0.0180786
R12988 iovss.n3100 iovss.n3099 0.0180786
R12989 iovss.n1103 iovss.n988 0.0180786
R12990 iovss.n1102 iovss.n987 0.0180786
R12991 iovss.n991 iovss.n990 0.0180786
R12992 iovss.n1035 iovss.n986 0.0180786
R12993 iovss.n993 iovss.n992 0.0180786
R12994 iovss.n1036 iovss.n985 0.0180786
R12995 iovss.n995 iovss.n994 0.0180786
R12996 iovss.n1037 iovss.n984 0.0180786
R12997 iovss.n997 iovss.n996 0.0180786
R12998 iovss.n1038 iovss.n983 0.0180786
R12999 iovss.n999 iovss.n998 0.0180786
R13000 iovss.n1039 iovss.n982 0.0180786
R13001 iovss.n1001 iovss.n1000 0.0180786
R13002 iovss.n1040 iovss.n981 0.0180786
R13003 iovss.n1003 iovss.n1002 0.0180786
R13004 iovss.n1041 iovss.n980 0.0180786
R13005 iovss.n1005 iovss.n1004 0.0180786
R13006 iovss.n1042 iovss.n979 0.0180786
R13007 iovss.n1007 iovss.n1006 0.0180786
R13008 iovss.n1043 iovss.n978 0.0180786
R13009 iovss.n1009 iovss.n1008 0.0180786
R13010 iovss.n1044 iovss.n977 0.0180786
R13011 iovss.n1011 iovss.n1010 0.0180786
R13012 iovss.n1045 iovss.n976 0.0180786
R13013 iovss.n1013 iovss.n1012 0.0180786
R13014 iovss.n1046 iovss.n975 0.0180786
R13015 iovss.n1015 iovss.n1014 0.0180786
R13016 iovss.n1047 iovss.n974 0.0180786
R13017 iovss.n1017 iovss.n1016 0.0180786
R13018 iovss.n1048 iovss.n973 0.0180786
R13019 iovss.n1019 iovss.n1018 0.0180786
R13020 iovss.n1049 iovss.n972 0.0180786
R13021 iovss.n1021 iovss.n1020 0.0180786
R13022 iovss.n1050 iovss.n971 0.0180786
R13023 iovss.n1023 iovss.n1022 0.0180786
R13024 iovss.n1051 iovss.n970 0.0180786
R13025 iovss.n1025 iovss.n1024 0.0180786
R13026 iovss.n1052 iovss.n969 0.0180786
R13027 iovss.n1027 iovss.n1026 0.0180786
R13028 iovss.n1053 iovss.n968 0.0180786
R13029 iovss.n1029 iovss.n1028 0.0180786
R13030 iovss.n1054 iovss.n967 0.0180786
R13031 iovss.n1031 iovss.n1030 0.0180786
R13032 iovss.n1055 iovss.n966 0.0180786
R13033 iovss.n1033 iovss.n1032 0.0180786
R13034 iovss.n3110 iovss.n963 0.0180786
R13035 iovss.n3112 iovss.n3111 0.0180786
R13036 iovss.n2764 iovss.n1318 0.0180786
R13037 iovss.n2768 iovss.n1318 0.0180786
R13038 iovss.n2766 iovss.n1316 0.0180786
R13039 iovss.n2771 iovss.n1316 0.0180786
R13040 iovss.n2774 iovss.n1313 0.0180786
R13041 iovss.n2775 iovss.n2774 0.0180786
R13042 iovss.n2790 iovss.n2789 0.0180786
R13043 iovss.n2789 iovss.n1226 0.0180786
R13044 iovss.n2795 iovss.n2792 0.0180786
R13045 iovss.n2792 iovss.n1227 0.0180786
R13046 iovss.n2800 iovss.n2797 0.0180786
R13047 iovss.n2797 iovss.n1228 0.0180786
R13048 iovss.n2805 iovss.n2802 0.0180786
R13049 iovss.n2802 iovss.n1229 0.0180786
R13050 iovss.n2810 iovss.n2807 0.0180786
R13051 iovss.n2807 iovss.n1230 0.0180786
R13052 iovss.n2815 iovss.n2812 0.0180786
R13053 iovss.n2812 iovss.n1231 0.0180786
R13054 iovss.n2820 iovss.n2817 0.0180786
R13055 iovss.n2817 iovss.n1232 0.0180786
R13056 iovss.n2825 iovss.n2822 0.0180786
R13057 iovss.n2822 iovss.n1233 0.0180786
R13058 iovss.n2830 iovss.n2827 0.0180786
R13059 iovss.n2827 iovss.n1234 0.0180786
R13060 iovss.n2835 iovss.n2832 0.0180786
R13061 iovss.n2832 iovss.n1235 0.0180786
R13062 iovss.n2840 iovss.n2837 0.0180786
R13063 iovss.n2837 iovss.n1236 0.0180786
R13064 iovss.n2845 iovss.n2842 0.0180786
R13065 iovss.n2842 iovss.n1237 0.0180786
R13066 iovss.n2850 iovss.n2847 0.0180786
R13067 iovss.n2847 iovss.n1238 0.0180786
R13068 iovss.n2855 iovss.n2852 0.0180786
R13069 iovss.n2852 iovss.n1239 0.0180786
R13070 iovss.n2860 iovss.n2857 0.0180786
R13071 iovss.n2857 iovss.n1240 0.0180786
R13072 iovss.n2865 iovss.n2862 0.0180786
R13073 iovss.n2862 iovss.n1241 0.0180786
R13074 iovss.n2870 iovss.n2867 0.0180786
R13075 iovss.n2867 iovss.n1242 0.0180786
R13076 iovss.n2875 iovss.n2872 0.0180786
R13077 iovss.n2872 iovss.n1243 0.0180786
R13078 iovss.n2880 iovss.n2877 0.0180786
R13079 iovss.n2877 iovss.n1244 0.0180786
R13080 iovss.n2885 iovss.n2882 0.0180786
R13081 iovss.n2882 iovss.n1245 0.0180786
R13082 iovss.n2889 iovss.n2888 0.0180786
R13083 iovss.n2889 iovss.n1246 0.0180786
R13084 iovss.n2899 iovss.n1247 0.0180786
R13085 iovss.n2899 iovss.n2898 0.0180786
R13086 iovss.n2790 iovss.n1225 0.0180786
R13087 iovss.n2794 iovss.n1226 0.0180786
R13088 iovss.n2795 iovss.n2794 0.0180786
R13089 iovss.n2799 iovss.n1227 0.0180786
R13090 iovss.n2800 iovss.n2799 0.0180786
R13091 iovss.n2804 iovss.n1228 0.0180786
R13092 iovss.n2805 iovss.n2804 0.0180786
R13093 iovss.n2809 iovss.n1229 0.0180786
R13094 iovss.n2810 iovss.n2809 0.0180786
R13095 iovss.n2814 iovss.n1230 0.0180786
R13096 iovss.n2815 iovss.n2814 0.0180786
R13097 iovss.n2819 iovss.n1231 0.0180786
R13098 iovss.n2820 iovss.n2819 0.0180786
R13099 iovss.n2824 iovss.n1232 0.0180786
R13100 iovss.n2825 iovss.n2824 0.0180786
R13101 iovss.n2829 iovss.n1233 0.0180786
R13102 iovss.n2830 iovss.n2829 0.0180786
R13103 iovss.n2834 iovss.n1234 0.0180786
R13104 iovss.n2835 iovss.n2834 0.0180786
R13105 iovss.n2839 iovss.n1235 0.0180786
R13106 iovss.n2840 iovss.n2839 0.0180786
R13107 iovss.n2844 iovss.n1236 0.0180786
R13108 iovss.n2845 iovss.n2844 0.0180786
R13109 iovss.n2849 iovss.n1237 0.0180786
R13110 iovss.n2850 iovss.n2849 0.0180786
R13111 iovss.n2854 iovss.n1238 0.0180786
R13112 iovss.n2855 iovss.n2854 0.0180786
R13113 iovss.n2859 iovss.n1239 0.0180786
R13114 iovss.n2860 iovss.n2859 0.0180786
R13115 iovss.n2864 iovss.n1240 0.0180786
R13116 iovss.n2865 iovss.n2864 0.0180786
R13117 iovss.n2869 iovss.n1241 0.0180786
R13118 iovss.n2870 iovss.n2869 0.0180786
R13119 iovss.n2874 iovss.n1242 0.0180786
R13120 iovss.n2875 iovss.n2874 0.0180786
R13121 iovss.n2879 iovss.n1243 0.0180786
R13122 iovss.n2880 iovss.n2879 0.0180786
R13123 iovss.n2884 iovss.n1244 0.0180786
R13124 iovss.n2885 iovss.n2884 0.0180786
R13125 iovss.n2887 iovss.n1245 0.0180786
R13126 iovss.n2888 iovss.n2887 0.0180786
R13127 iovss.n2892 iovss.n1246 0.0180786
R13128 iovss.n2892 iovss.n1247 0.0180786
R13129 iovss.n2898 iovss.n2897 0.0180786
R13130 iovss.n1342 iovss.n1338 0.0180786
R13131 iovss.n2759 iovss.n1347 0.0180786
R13132 iovss.n1348 iovss.n1343 0.0180786
R13133 iovss.n1346 iovss.n1345 0.0180786
R13134 iovss.n1381 iovss.n1380 0.0180786
R13135 iovss.n2718 iovss.n1344 0.0180786
R13136 iovss.n2710 iovss.n2604 0.0180786
R13137 iovss.n2750 iovss.n2708 0.0180786
R13138 iovss.n2707 iovss.n2606 0.0180786
R13139 iovss.n2749 iovss.n2705 0.0180786
R13140 iovss.n2704 iovss.n2608 0.0180786
R13141 iovss.n2748 iovss.n2702 0.0180786
R13142 iovss.n2701 iovss.n2610 0.0180786
R13143 iovss.n2747 iovss.n2699 0.0180786
R13144 iovss.n2698 iovss.n2612 0.0180786
R13145 iovss.n2746 iovss.n2696 0.0180786
R13146 iovss.n2695 iovss.n2614 0.0180786
R13147 iovss.n2745 iovss.n2693 0.0180786
R13148 iovss.n2692 iovss.n2616 0.0180786
R13149 iovss.n2744 iovss.n2690 0.0180786
R13150 iovss.n2689 iovss.n2618 0.0180786
R13151 iovss.n2743 iovss.n2687 0.0180786
R13152 iovss.n2686 iovss.n2620 0.0180786
R13153 iovss.n2742 iovss.n2684 0.0180786
R13154 iovss.n2683 iovss.n2622 0.0180786
R13155 iovss.n2741 iovss.n2681 0.0180786
R13156 iovss.n2680 iovss.n2624 0.0180786
R13157 iovss.n2740 iovss.n2678 0.0180786
R13158 iovss.n2677 iovss.n2626 0.0180786
R13159 iovss.n2739 iovss.n2675 0.0180786
R13160 iovss.n2674 iovss.n2628 0.0180786
R13161 iovss.n2738 iovss.n2672 0.0180786
R13162 iovss.n2671 iovss.n2630 0.0180786
R13163 iovss.n2737 iovss.n2669 0.0180786
R13164 iovss.n2668 iovss.n2632 0.0180786
R13165 iovss.n2736 iovss.n2666 0.0180786
R13166 iovss.n2665 iovss.n2634 0.0180786
R13167 iovss.n2735 iovss.n2663 0.0180786
R13168 iovss.n2662 iovss.n2636 0.0180786
R13169 iovss.n2734 iovss.n2660 0.0180786
R13170 iovss.n2659 iovss.n2638 0.0180786
R13171 iovss.n2733 iovss.n2657 0.0180786
R13172 iovss.n2656 iovss.n2640 0.0180786
R13173 iovss.n2732 iovss.n2654 0.0180786
R13174 iovss.n2653 iovss.n2642 0.0180786
R13175 iovss.n2731 iovss.n2651 0.0180786
R13176 iovss.n2650 iovss.n2644 0.0180786
R13177 iovss.n2730 iovss.n2648 0.0180786
R13178 iovss.n2647 iovss.n2645 0.0180786
R13179 iovss.n2754 iovss.n1409 0.0180786
R13180 iovss.n2645 iovss.n1409 0.0180786
R13181 iovss.n2648 iovss.n2647 0.0180786
R13182 iovss.n2730 iovss.n2644 0.0180786
R13183 iovss.n2651 iovss.n2650 0.0180786
R13184 iovss.n2731 iovss.n2642 0.0180786
R13185 iovss.n2654 iovss.n2653 0.0180786
R13186 iovss.n2732 iovss.n2640 0.0180786
R13187 iovss.n2657 iovss.n2656 0.0180786
R13188 iovss.n2733 iovss.n2638 0.0180786
R13189 iovss.n2660 iovss.n2659 0.0180786
R13190 iovss.n2734 iovss.n2636 0.0180786
R13191 iovss.n2663 iovss.n2662 0.0180786
R13192 iovss.n2735 iovss.n2634 0.0180786
R13193 iovss.n2666 iovss.n2665 0.0180786
R13194 iovss.n2736 iovss.n2632 0.0180786
R13195 iovss.n2669 iovss.n2668 0.0180786
R13196 iovss.n2737 iovss.n2630 0.0180786
R13197 iovss.n2672 iovss.n2671 0.0180786
R13198 iovss.n2738 iovss.n2628 0.0180786
R13199 iovss.n2675 iovss.n2674 0.0180786
R13200 iovss.n2739 iovss.n2626 0.0180786
R13201 iovss.n2678 iovss.n2677 0.0180786
R13202 iovss.n2740 iovss.n2624 0.0180786
R13203 iovss.n2681 iovss.n2680 0.0180786
R13204 iovss.n2741 iovss.n2622 0.0180786
R13205 iovss.n2684 iovss.n2683 0.0180786
R13206 iovss.n2742 iovss.n2620 0.0180786
R13207 iovss.n2687 iovss.n2686 0.0180786
R13208 iovss.n2743 iovss.n2618 0.0180786
R13209 iovss.n2690 iovss.n2689 0.0180786
R13210 iovss.n2744 iovss.n2616 0.0180786
R13211 iovss.n2693 iovss.n2692 0.0180786
R13212 iovss.n2745 iovss.n2614 0.0180786
R13213 iovss.n2696 iovss.n2695 0.0180786
R13214 iovss.n2746 iovss.n2612 0.0180786
R13215 iovss.n2699 iovss.n2698 0.0180786
R13216 iovss.n2747 iovss.n2610 0.0180786
R13217 iovss.n2702 iovss.n2701 0.0180786
R13218 iovss.n2748 iovss.n2608 0.0180786
R13219 iovss.n2705 iovss.n2704 0.0180786
R13220 iovss.n2749 iovss.n2606 0.0180786
R13221 iovss.n2708 iovss.n2707 0.0180786
R13222 iovss.n2750 iovss.n2604 0.0180786
R13223 iovss.n2711 iovss.n2710 0.0180786
R13224 iovss.n1381 iovss.n1344 0.0180786
R13225 iovss.n1380 iovss.n1346 0.0180786
R13226 iovss.n1345 iovss.n1343 0.0180786
R13227 iovss.n2759 iovss.n1348 0.0180786
R13228 iovss.n1347 iovss.n1342 0.0180786
R13229 iovss.n2761 iovss.n1338 0.0180786
R13230 iovss.n2765 iovss.n2764 0.0180786
R13231 iovss.n2769 iovss.n2768 0.0180786
R13232 iovss.n2769 iovss.n2766 0.0180786
R13233 iovss.n2772 iovss.n2771 0.0180786
R13234 iovss.n2772 iovss.n1313 0.0180786
R13235 iovss.n2776 iovss.n2775 0.0180786
R13236 iovss.n894 iovss.n893 0.0180786
R13237 iovss.n3139 iovss.n891 0.0180786
R13238 iovss.n896 iovss.n895 0.0180786
R13239 iovss.n3140 iovss.n890 0.0180786
R13240 iovss.n898 iovss.n897 0.0180786
R13241 iovss.n3141 iovss.n889 0.0180786
R13242 iovss.n900 iovss.n899 0.0180786
R13243 iovss.n3142 iovss.n888 0.0180786
R13244 iovss.n902 iovss.n901 0.0180786
R13245 iovss.n3143 iovss.n887 0.0180786
R13246 iovss.n3145 iovss.n903 0.0180786
R13247 iovss.n1196 iovss.n915 0.0180786
R13248 iovss.n917 iovss.n916 0.0180786
R13249 iovss.n1197 iovss.n911 0.0180786
R13250 iovss.n922 iovss.n921 0.0180786
R13251 iovss.n1195 iovss.n924 0.0180786
R13252 iovss.n3135 iovss.n926 0.0180786
R13253 iovss.n925 iovss.n908 0.0180786
R13254 iovss.n3137 iovss.n906 0.0180786
R13255 iovss.n940 iovss.n939 0.0180786
R13256 iovss.n946 iovss.n937 0.0180786
R13257 iovss.n942 iovss.n941 0.0180786
R13258 iovss.n947 iovss.n936 0.0180786
R13259 iovss.n944 iovss.n943 0.0180786
R13260 iovss.n948 iovss.n935 0.0180786
R13261 iovss.n3129 iovss.n951 0.0180786
R13262 iovss.n950 iovss.n934 0.0180786
R13263 iovss.n3131 iovss.n929 0.0180786
R13264 iovss.n933 iovss.n928 0.0180786
R13265 iovss.n931 iovss.n905 0.0180786
R13266 iovss.n1174 iovss.n1124 0.0180349
R13267 iovss.n1213 iovss.n1164 0.0180327
R13268 iovss.n918 iovss.n917 0.0180322
R13269 iovss.n1147 iovss.n1146 0.0180322
R13270 iovss.n1209 iovss.n1184 0.0180322
R13271 iovss.n1207 iovss.n1191 0.0180306
R13272 iovss.n1154 iovss.n1132 0.0180294
R13273 iovss.n1208 iovss.n1117 0.0180294
R13274 iovss.n3086 iovss.n1130 0.0180294
R13275 iovss.n1217 iovss.n1144 0.0180284
R13276 iovss.n1181 iovss.n1180 0.0180266
R13277 iovss.n1167 iovss.n1166 0.0180266
R13278 iovss.n920 iovss.n910 0.0180266
R13279 iovss.n3090 iovss.n1122 0.0180239
R13280 iovss.n1172 iovss.n1125 0.0180239
R13281 iovss.n1203 iovss.n1202 0.0180219
R13282 iovss.n1187 iovss.n1186 0.0180211
R13283 iovss.n1161 iovss.n1160 0.0180211
R13284 iovss.n1150 iovss.n1149 0.0180211
R13285 iovss.n1189 iovss.n1118 0.0180184
R13286 iovss.n1156 iovss.n1129 0.0180184
R13287 iovss.n1152 iovss.n1133 0.0180184
R13288 iovss.n923 iovss.n909 0.0180156
R13289 iovss.n1141 iovss.n1140 0.0180156
R13290 iovss.n1178 iovss.n1176 0.0180156
R13291 iovss.n1170 iovss.n1169 0.0180156
R13292 iovss.n1193 iovss.n913 0.0180153
R13293 iovss.n1194 iovss.n1193 0.0180132
R13294 iovss.n1176 iovss.n1121 0.0180129
R13295 iovss.n1169 iovss.n1126 0.0180129
R13296 iovss.n924 iovss.n923 0.0180129
R13297 iovss.n1140 iovss.n1136 0.0180129
R13298 iovss.n1153 iovss.n1152 0.0180101
R13299 iovss.n1190 iovss.n1189 0.0180101
R13300 iovss.n1158 iovss.n1156 0.0180101
R13301 iovss.n1149 iovss.n1134 0.0180073
R13302 iovss.n1186 iovss.n1119 0.0180073
R13303 iovss.n1160 iovss.n1128 0.0180073
R13304 iovss.n1202 iovss.n1201 0.0180066
R13305 iovss.n3091 iovss.n3090 0.0180046
R13306 iovss.n1173 iovss.n1172 0.0180046
R13307 iovss.n922 iovss.n920 0.0180018
R13308 iovss.n1180 iovss.n1120 0.0180018
R13309 iovss.n1166 iovss.n1127 0.0180018
R13310 iovss.n1218 iovss.n1217 0.018
R13311 iovss.n3096 iovss.n1208 0.017999
R13312 iovss.n3087 iovss.n3086 0.017999
R13313 iovss.n1155 iovss.n1154 0.017999
R13314 iovss.n1204 iovss.n1191 0.0179979
R13315 iovss.n1210 iovss.n1209 0.0179962
R13316 iovss.n919 iovss.n918 0.0179962
R13317 iovss.n1146 iovss.n1135 0.0179962
R13318 iovss.n1214 iovss.n1213 0.0179957
R13319 iovss.n1175 iovss.n1174 0.0179935
R13320 iovss.n1379 iovss.n1378 0.0179603
R13321 iovss.n2700 iovss.n1371 0.0179603
R13322 iovss.n2670 iovss.n1360 0.0179603
R13323 iovss.n2649 iovss.n1405 0.0179603
R13324 iovss.n2770 iovss.n1279 0.0179603
R13325 iovss.n2803 iovss.n1269 0.0179603
R13326 iovss.n2853 iovss.n1258 0.0179603
R13327 iovss.n1304 iovss.n1303 0.0179603
R13328 iovss.n2725 iovss.n1385 0.0175485
R13329 iovss.n2709 iovss.n1387 0.0175485
R13330 iovss.n2661 iovss.n1357 0.0175485
R13331 iovss.n2658 iovss.n1355 0.0175485
R13332 iovss.n2783 iovss.n1282 0.0175485
R13333 iovss.n1285 iovss.n1284 0.0175485
R13334 iovss.n2868 iovss.n1255 0.0175485
R13335 iovss.n2873 iovss.n1253 0.0175485
R13336 iovss.n2617 iovss.n1393 0.0170873
R13337 iovss.n2619 iovss.n1394 0.0170873
R13338 iovss.n2821 iovss.n1291 0.0170873
R13339 iovss.n2826 iovss.n1292 0.0170873
R13340 iovss.n1377 iovss.n1351 0.0166755
R13341 iovss.n2609 iovss.n1370 0.0166755
R13342 iovss.n2627 iovss.n1399 0.0166755
R13343 iovss.n2643 iovss.n1406 0.0166755
R13344 iovss.n1315 iovss.n1275 0.0166755
R13345 iovss.n2801 iovss.n1268 0.0166755
R13346 iovss.n2846 iovss.n1297 0.0166755
R13347 iovss.n2891 iovss.n2890 0.0166755
R13348 iovss.n2685 iovss.n1364 0.0165499
R13349 iovss.n2828 iovss.n1262 0.0165499
R13350 iovss.n2758 iovss.n1350 0.0162143
R13351 iovss.n2697 iovss.n1369 0.0162143
R13352 iovss.n2673 iovss.n1361 0.0162143
R13353 iovss.n2646 iovss.n1407 0.0162143
R13354 iovss.n2767 iovss.n1278 0.0162143
R13355 iovss.n2808 iovss.n1267 0.0162143
R13356 iovss.n2848 iovss.n1259 0.0162143
R13357 iovss.n2894 iovss.n2893 0.0162143
R13358 iovss.n2727 iovss.n1374 0.0153413
R13359 iovss.n2727 iovss.n1386 0.0153413
R13360 iovss.n2635 iovss.n1402 0.0153413
R13361 iovss.n2635 iovss.n1356 0.0153413
R13362 iovss.n2755 iovss 0.0153413
R13363 iovss.n2785 iovss.n1272 0.0153413
R13364 iovss.n2785 iovss.n1283 0.0153413
R13365 iovss.n2866 iovss.n1300 0.0153413
R13366 iovss.n2866 iovss.n1254 0.0153413
R13367 iovss.n2896 iovss 0.0153413
R13368 iovss.n2092 iovss.n1996 0.0148733
R13369 iovss.n2562 iovss.n1485 0.0148733
R13370 iovss.n2452 iovss.n1439 0.0148733
R13371 iovss.n2567 iovss.n1439 0.0148733
R13372 iovss.n2568 iovss.n2567 0.0148733
R13373 iovss.n2569 iovss.n2568 0.0148733
R13374 iovss.n2573 iovss.n2572 0.0148733
R13375 iovss.n2574 iovss.n2573 0.0148733
R13376 iovss.n2574 iovss.n1434 0.0148733
R13377 iovss.n2586 iovss.n1435 0.0148733
R13378 iovss.n2582 iovss.n1435 0.0148733
R13379 iovss.n2582 iovss.n2581 0.0148733
R13380 iovss.n2579 iovss.n1412 0.0148733
R13381 iovss.n2599 iovss.n1412 0.0148733
R13382 iovss.n2599 iovss.n2598 0.0148733
R13383 iovss.n1419 iovss.n1413 0.0148733
R13384 iovss.n1420 iovss.n1419 0.0148733
R13385 iovss.n1420 iovss.n1415 0.0148733
R13386 iovss.n1424 iovss.n1416 0.0148733
R13387 iovss.n2566 iovss.n2565 0.0148733
R13388 iovss.n2566 iovss.n1438 0.0148733
R13389 iovss.n2570 iovss.n1438 0.0148733
R13390 iovss.n2571 iovss.n2570 0.0148733
R13391 iovss.n2571 iovss.n1436 0.0148733
R13392 iovss.n2575 iovss.n1436 0.0148733
R13393 iovss.n2576 iovss.n2575 0.0148733
R13394 iovss.n2585 iovss.n2576 0.0148733
R13395 iovss.n2585 iovss.n2584 0.0148733
R13396 iovss.n2584 iovss.n2583 0.0148733
R13397 iovss.n2583 iovss.n2577 0.0148733
R13398 iovss.n2578 iovss.n2577 0.0148733
R13399 iovss.n2578 iovss.n1410 0.0148733
R13400 iovss.n2600 iovss.n1411 0.0148733
R13401 iovss.n1417 iovss.n1411 0.0148733
R13402 iovss.n1418 iovss.n1417 0.0148733
R13403 iovss.n1421 iovss.n1418 0.0148733
R13404 iovss.n1422 iovss.n1421 0.0148733
R13405 iovss.n1423 iovss.n1422 0.0148733
R13406 iovss.n1423 iovss.n1249 0.0148733
R13407 iovss.n2063 iovss.n2009 0.01458
R13408 iovss.n2454 iovss.n2453 0.01458
R13409 iovss.n2758 iovss.n2757 0.0144683
R13410 iovss.n2697 iovss.n1390 0.0144683
R13411 iovss.n2673 iovss.n1398 0.0144683
R13412 iovss.n2646 iovss.n1352 0.0144683
R13413 iovss.n2767 iovss.n1276 0.0144683
R13414 iovss.n2808 iovss.n1288 0.0144683
R13415 iovss.n2848 iovss.n1296 0.0144683
R13416 iovss.n2893 iovss.n1250 0.0144683
R13417 iovss.n2065 iovss.n2006 0.0139933
R13418 iovss.n2572 iovss.n1437 0.0139933
R13419 iovss.n2521 iovss.n1474 0.0137
R13420 iovss.n2518 iovss.n1469 0.0137
R13421 iovss.n2617 iovss.n1365 0.0135952
R13422 iovss.n2821 iovss.n1263 0.0135952
R13423 iovss.n2043 iovss.n2011 0.0134067
R13424 iovss.n2461 iovss.n2451 0.0134067
R13425 iovss.n2067 iovss.n2004 0.01282
R13426 iovss.n2587 iovss.n2586 0.01282
R13427 iovss.n2931 iovss 0.0127222
R13428 iovss.n1514 iovss.n1476 0.0125267
R13429 iovss.n1545 iovss.n1537 0.0125267
R13430 iovss.n2072 iovss.n2071 0.0125
R13431 iovss.n2071 iovss.n2070 0.0125
R13432 iovss.n2070 iovss.n2041 0.0125
R13433 iovss.n2061 iovss.n2041 0.0125
R13434 iovss.n2061 iovss.n2060 0.0125
R13435 iovss.n2060 iovss.n2059 0.0125
R13436 iovss.n2059 iovss.n2052 0.0125
R13437 iovss.n2052 iovss.n1508 0.0125
R13438 iovss.n2537 iovss.n1508 0.0125
R13439 iovss.n2537 iovss.n2536 0.0125
R13440 iovss.n2536 iovss.n2535 0.0125
R13441 iovss.n2535 iovss.n1512 0.0125
R13442 iovss.n2526 iovss.n1512 0.0125
R13443 iovss.n2526 iovss.n2525 0.0125
R13444 iovss.n2525 iovss.n2524 0.0125
R13445 iovss.n2524 iovss.n1521 0.0125
R13446 iovss.n2516 iovss.n1521 0.0125
R13447 iovss.n2516 iovss.n2515 0.0125
R13448 iovss.n2515 iovss.n2514 0.0125
R13449 iovss.n2514 iovss.n1529 0.0125
R13450 iovss.n2490 iovss.n1529 0.0125
R13451 iovss.n2490 iovss.n2489 0.0125
R13452 iovss.n2489 iovss.n2488 0.0125
R13453 iovss.n2488 iovss.n2410 0.0125
R13454 iovss.n2466 iovss.n2410 0.0125
R13455 iovss.n2466 iovss.n2465 0.0125
R13456 iovss.n2465 iovss.n2464 0.0125
R13457 iovss.n2464 iovss.n2435 0.0125
R13458 iovss.n2435 iovss.n1431 0.0125
R13459 iovss.n2590 iovss.n1431 0.0125
R13460 iovss.n2590 iovss.n1429 0.0125
R13461 iovss.n2594 iovss.n1429 0.0125
R13462 iovss.n3250 iovss.n673 0.0124589
R13463 iovss.n3393 iovss.n303 0.0124589
R13464 iovss.n3428 iovss.n220 0.0124589
R13465 iovss.n2056 iovss.n2013 0.0122333
R13466 iovss.n2444 iovss.n2443 0.0122333
R13467 iovss.n2601 iovss.n2600 0.0122333
R13468 iovss.n579 iovss.n578 0.0119199
R13469 iovss.n1539 iovss.n1535 0.0117671
R13470 iovss.n1544 iovss.n1543 0.0117671
R13471 iovss.n1546 iovss.n1535 0.0117671
R13472 iovss.n1543 iovss.n1538 0.0117671
R13473 iovss.n1534 iovss.n1442 0.0117671
R13474 iovss.n1538 iovss.n1533 0.0117671
R13475 iovss.n1539 iovss.n1534 0.0117671
R13476 iovss.n1533 iovss.n1445 0.0117671
R13477 iovss.n1990 iovss.n1987 0.0117136
R13478 iovss.n1986 iovss.n1446 0.0117136
R13479 iovss.n1989 iovss.n1983 0.0117136
R13480 iovss.n1995 iovss.n1988 0.0117136
R13481 iovss.n1990 iovss.n1984 0.0117136
R13482 iovss.n1987 iovss.n1986 0.0117136
R13483 iovss.n1989 iovss.n1447 0.0117136
R13484 iovss.n1988 iovss.n1983 0.0117136
R13485 iovss.n2035 iovss.n2002 0.0116467
R13486 iovss.n2580 iovss.n2579 0.0116467
R13487 iovss.n694 iovss.n334 0.0116063
R13488 iovss.n3413 iovss.n3395 0.0115591
R13489 iovss.n577 iovss.n576 0.0115
R13490 iovss.n576 iovss.n575 0.0115
R13491 iovss.n575 iovss.n573 0.0115
R13492 iovss.n585 iovss.n573 0.0115
R13493 iovss.n585 iovss.n584 0.0115
R13494 iovss.n584 iovss.n574 0.0115
R13495 iovss.n574 iovss.n569 0.0115
R13496 iovss.n591 iovss.n569 0.0115
R13497 iovss.n592 iovss.n591 0.0115
R13498 iovss.n592 iovss.n566 0.0115
R13499 iovss.n597 iovss.n566 0.0115
R13500 iovss.n599 iovss.n597 0.0115
R13501 iovss.n599 iovss.n598 0.0115
R13502 iovss.n598 iovss.n560 0.0115
R13503 iovss.n606 iovss.n560 0.0115
R13504 iovss.n606 iovss.n605 0.0115
R13505 iovss.n605 iovss.n562 0.0115
R13506 iovss.n562 iovss.n561 0.0115
R13507 iovss.n561 iovss.n486 0.0115
R13508 iovss.n3264 iovss.n486 0.0115
R13509 iovss.n3264 iovss.n3263 0.0115
R13510 iovss.n3263 iovss.n487 0.0115
R13511 iovss.n487 iovss.n482 0.0115
R13512 iovss.n3270 iovss.n482 0.0115
R13513 iovss.n3272 iovss.n3270 0.0115
R13514 iovss.n3272 iovss.n3271 0.0115
R13515 iovss.n3271 iovss.n479 0.0115
R13516 iovss.n3280 iovss.n479 0.0115
R13517 iovss.n3280 iovss.n3279 0.0115
R13518 iovss.n3279 iovss.n480 0.0115
R13519 iovss.n480 iovss.n475 0.0115
R13520 iovss.n3286 iovss.n475 0.0115
R13521 iovss.n3287 iovss.n3286 0.0115
R13522 iovss.n3287 iovss.n472 0.0115
R13523 iovss.n3292 iovss.n472 0.0115
R13524 iovss.n3295 iovss.n3292 0.0115
R13525 iovss.n3295 iovss.n3294 0.0115
R13526 iovss.n3294 iovss.n3293 0.0115
R13527 iovss.n3293 iovss.n454 0.0115
R13528 iovss.n3300 iovss.n454 0.0115
R13529 iovss.n3300 iovss.n455 0.0115
R13530 iovss.n3302 iovss.n455 0.0115
R13531 iovss.n3302 iovss.n456 0.0115
R13532 iovss.n3304 iovss.n456 0.0115
R13533 iovss.n3304 iovss.n457 0.0115
R13534 iovss.n466 iovss.n457 0.0115
R13535 iovss.n466 iovss.n458 0.0115
R13536 iovss.n3309 iovss.n458 0.0115
R13537 iovss.n3309 iovss.n459 0.0115
R13538 iovss.n3311 iovss.n459 0.0115
R13539 iovss.n3311 iovss.n460 0.0115
R13540 iovss.n3313 iovss.n460 0.0115
R13541 iovss.n3313 iovss.n461 0.0115
R13542 iovss.n462 iovss.n461 0.0115
R13543 iovss.n3320 iovss.n462 0.0115
R13544 iovss.n3320 iovss.n3319 0.0115
R13545 iovss.n3319 iovss.n463 0.0115
R13546 iovss.n463 iovss.n76 0.0115
R13547 iovss.n3439 iovss.n76 0.0115
R13548 iovss.n3441 iovss.n3439 0.0115
R13549 iovss.n3441 iovss.n3440 0.0115
R13550 iovss.n3440 iovss.n70 0.0115
R13551 iovss.n3449 iovss.n70 0.0115
R13552 iovss.n3449 iovss.n3448 0.0115
R13553 iovss.n3448 iovss.n71 0.0115
R13554 iovss.n71 iovss.n66 0.0115
R13555 iovss.n3455 iovss.n66 0.0115
R13556 iovss.n3456 iovss.n3455 0.0115
R13557 iovss.n3457 iovss.n3456 0.0115
R13558 iovss.n3458 iovss.n3457 0.0115
R13559 iovss.n3458 iovss.n60 0.0115
R13560 iovss.n62 iovss.n60 0.0115
R13561 iovss.n62 iovss.n61 0.0115
R13562 iovss.n3464 iovss.n61 0.0115
R13563 iovss.n2528 iovss.n1478 0.0113533
R13564 iovss.n2511 iovss.n2510 0.0113533
R13565 iovss.n2564 iovss.n1442 0.01128
R13566 iovss.n2564 iovss.n1445 0.01128
R13567 iovss.n2564 iovss.n1446 0.0112264
R13568 iovss.n2564 iovss.n1447 0.0112264
R13569 iovss.n2054 iovss.n2015 0.01106
R13570 iovss.n2470 iovss.n2469 0.01106
R13571 iovss.n2074 iovss.n2000 0.0104733
R13572 iovss.n2597 iovss.n1413 0.0104733
R13573 iovss.n2530 iovss.n1480 0.01018
R13574 iovss.n2501 iovss.n2500 0.01018
R13575 iovss.n1991 iovss.n1985 0.00988667
R13576 iovss.n2478 iovss.n2477 0.00988667
R13577 iovss.n2077 iovss.n1999 0.0093
R13578 iovss.n1425 iovss.n1424 0.0093
R13579 iovss.n2532 iovss.n1482 0.00900667
R13580 iovss.n2493 iovss.n2403 0.00900667
R13581 iovss.n2558 iovss.n2540 0.00871333
R13582 iovss.n2485 iovss.n2426 0.00871333
R13583 iovss.n614 iovss.n380 0.0082
R13584 iovss.n2090 iovss.n1962 0.00818093
R13585 iovss.n2078 iovss.n1963 0.00818093
R13586 iovss.n2081 iovss.n2080 0.00818093
R13587 iovss.n2033 iovss.n1964 0.00818093
R13588 iovss.n2032 iovss.n1965 0.00818093
R13589 iovss.n2082 iovss.n2001 0.00818093
R13590 iovss.n2031 iovss.n1966 0.00818093
R13591 iovss.n2030 iovss.n1967 0.00818093
R13592 iovss.n2083 iovss.n2003 0.00818093
R13593 iovss.n2029 iovss.n1968 0.00818093
R13594 iovss.n2028 iovss.n1969 0.00818093
R13595 iovss.n2084 iovss.n2005 0.00818093
R13596 iovss.n2027 iovss.n1970 0.00818093
R13597 iovss.n2026 iovss.n1971 0.00818093
R13598 iovss.n2085 iovss.n2007 0.00818093
R13599 iovss.n2025 iovss.n1972 0.00818093
R13600 iovss.n2023 iovss.n2008 0.00818093
R13601 iovss.n2009 iovss.n1974 0.00818093
R13602 iovss.n2086 iovss.n2010 0.00818093
R13603 iovss.n2010 iovss.n1975 0.00818093
R13604 iovss.n2011 iovss.n1976 0.00818093
R13605 iovss.n2087 iovss.n2012 0.00818093
R13606 iovss.n2012 iovss.n1977 0.00818093
R13607 iovss.n2013 iovss.n1978 0.00818093
R13608 iovss.n2088 iovss.n2014 0.00818093
R13609 iovss.n2014 iovss.n1979 0.00818093
R13610 iovss.n2015 iovss.n1980 0.00818093
R13611 iovss.n2092 iovss.n1981 0.00818093
R13612 iovss.n1992 iovss.n1991 0.00818093
R13613 iovss.n1993 iovss.n1485 0.00818093
R13614 iovss.n2559 iovss.n2558 0.00818093
R13615 iovss.n2555 iovss.n1450 0.00818093
R13616 iovss.n2555 iovss.n2554 0.00818093
R13617 iovss.n1487 iovss.n1451 0.00818093
R13618 iovss.n2541 iovss.n1452 0.00818093
R13619 iovss.n1488 iovss.n1452 0.00818093
R13620 iovss.n1489 iovss.n1453 0.00818093
R13621 iovss.n2542 iovss.n1454 0.00818093
R13622 iovss.n1490 iovss.n1454 0.00818093
R13623 iovss.n1491 iovss.n1455 0.00818093
R13624 iovss.n2543 iovss.n1456 0.00818093
R13625 iovss.n1492 iovss.n1456 0.00818093
R13626 iovss.n1493 iovss.n1457 0.00818093
R13627 iovss.n2544 iovss.n1458 0.00818093
R13628 iovss.n1494 iovss.n1458 0.00818093
R13629 iovss.n1495 iovss.n1459 0.00818093
R13630 iovss.n2545 iovss.n1460 0.00818093
R13631 iovss.n1496 iovss.n1460 0.00818093
R13632 iovss.n1497 iovss.n1461 0.00818093
R13633 iovss.n2546 iovss.n1462 0.00818093
R13634 iovss.n1498 iovss.n1462 0.00818093
R13635 iovss.n2547 iovss.n1463 0.00818093
R13636 iovss.n1499 iovss.n1463 0.00818093
R13637 iovss.n2548 iovss.n1464 0.00818093
R13638 iovss.n1500 iovss.n1464 0.00818093
R13639 iovss.n2549 iovss.n1465 0.00818093
R13640 iovss.n2550 iovss.n1466 0.00818093
R13641 iovss.n1501 iovss.n1466 0.00818093
R13642 iovss.n2551 iovss.n1467 0.00818093
R13643 iovss.n1542 iovss.n1540 0.00818093
R13644 iovss.n1542 iovss.n1541 0.00818093
R13645 iovss.n1547 iovss.n1532 0.00818093
R13646 iovss.n2509 iovss.n2508 0.00818093
R13647 iovss.n2508 iovss.n2506 0.00818093
R13648 iovss.n2504 iovss.n2503 0.00818093
R13649 iovss.n2499 iovss.n2498 0.00818093
R13650 iovss.n2498 iovss.n2497 0.00818093
R13651 iovss.n2495 iovss.n2494 0.00818093
R13652 iovss.n2414 iovss.n2413 0.00818093
R13653 iovss.n2415 iovss.n2414 0.00818093
R13654 iovss.n2418 iovss.n2417 0.00818093
R13655 iovss.n2422 iovss.n2421 0.00818093
R13656 iovss.n2423 iovss.n2422 0.00818093
R13657 iovss.n2426 iovss.n2425 0.00818093
R13658 iovss.n2483 iovss.n2482 0.00818093
R13659 iovss.n2482 iovss.n2481 0.00818093
R13660 iovss.n2479 iovss.n2478 0.00818093
R13661 iovss.n2475 iovss.n2474 0.00818093
R13662 iovss.n2474 iovss.n2473 0.00818093
R13663 iovss.n2471 iovss.n2470 0.00818093
R13664 iovss.n2439 iovss.n2438 0.00818093
R13665 iovss.n2440 iovss.n2439 0.00818093
R13666 iovss.n2443 iovss.n2442 0.00818093
R13667 iovss.n2447 iovss.n2446 0.00818093
R13668 iovss.n2448 iovss.n2447 0.00818093
R13669 iovss.n2451 iovss.n2450 0.00818093
R13670 iovss.n2459 iovss.n2458 0.00818093
R13671 iovss.n2458 iovss.n2457 0.00818093
R13672 iovss.n2455 iovss.n2454 0.00818093
R13673 iovss.n2016 iovss.n1980 0.00818093
R13674 iovss.n2017 iovss.n1979 0.00818093
R13675 iovss.n2018 iovss.n1978 0.00818093
R13676 iovss.n2019 iovss.n1977 0.00818093
R13677 iovss.n2020 iovss.n1976 0.00818093
R13678 iovss.n2021 iovss.n1975 0.00818093
R13679 iovss.n2022 iovss.n1974 0.00818093
R13680 iovss.n2008 iovss.n1972 0.00818093
R13681 iovss.n2007 iovss.n1971 0.00818093
R13682 iovss.n2006 iovss.n1970 0.00818093
R13683 iovss.n2005 iovss.n1969 0.00818093
R13684 iovss.n2004 iovss.n1968 0.00818093
R13685 iovss.n2003 iovss.n1967 0.00818093
R13686 iovss.n2002 iovss.n1966 0.00818093
R13687 iovss.n2001 iovss.n1965 0.00818093
R13688 iovss.n2000 iovss.n1964 0.00818093
R13689 iovss.n2080 iovss.n1963 0.00818093
R13690 iovss.n1999 iovss.n1962 0.00818093
R13691 iovss.n2016 iovss.n1981 0.00818093
R13692 iovss.n2088 iovss.n2018 0.00818093
R13693 iovss.n2087 iovss.n2020 0.00818093
R13694 iovss.n2086 iovss.n2022 0.00818093
R13695 iovss.n2085 iovss.n2025 0.00818093
R13696 iovss.n2084 iovss.n2027 0.00818093
R13697 iovss.n2083 iovss.n2029 0.00818093
R13698 iovss.n2082 iovss.n2031 0.00818093
R13699 iovss.n2081 iovss.n2033 0.00818093
R13700 iovss.n2024 iovss.n2023 0.00818093
R13701 iovss.n1541 iovss.n1536 0.00818093
R13702 iovss.n1545 iovss.n1540 0.00818093
R13703 iovss.n1536 iovss.n1532 0.00818093
R13704 iovss.n1994 iovss.n1993 0.00818093
R13705 iovss.n1994 iovss.n1992 0.00818093
R13706 iovss.n1501 iovss.n1468 0.00818093
R13707 iovss.n1500 iovss.n1470 0.00818093
R13708 iovss.n1499 iovss.n1471 0.00818093
R13709 iovss.n1498 iovss.n1472 0.00818093
R13710 iovss.n1497 iovss.n1473 0.00818093
R13711 iovss.n1496 iovss.n1474 0.00818093
R13712 iovss.n1495 iovss.n1475 0.00818093
R13713 iovss.n1494 iovss.n1476 0.00818093
R13714 iovss.n1493 iovss.n1477 0.00818093
R13715 iovss.n1492 iovss.n1478 0.00818093
R13716 iovss.n1491 iovss.n1479 0.00818093
R13717 iovss.n1490 iovss.n1480 0.00818093
R13718 iovss.n1489 iovss.n1481 0.00818093
R13719 iovss.n1488 iovss.n1482 0.00818093
R13720 iovss.n1487 iovss.n1483 0.00818093
R13721 iovss.n2554 iovss.n1484 0.00818093
R13722 iovss.n2551 iovss.n1468 0.00818093
R13723 iovss.n2550 iovss.n1469 0.00818093
R13724 iovss.n2549 iovss.n1470 0.00818093
R13725 iovss.n2548 iovss.n1471 0.00818093
R13726 iovss.n2547 iovss.n1472 0.00818093
R13727 iovss.n2546 iovss.n1473 0.00818093
R13728 iovss.n2545 iovss.n1475 0.00818093
R13729 iovss.n2544 iovss.n1477 0.00818093
R13730 iovss.n2543 iovss.n1479 0.00818093
R13731 iovss.n2542 iovss.n1481 0.00818093
R13732 iovss.n2541 iovss.n1483 0.00818093
R13733 iovss.n2560 iovss.n2559 0.00818093
R13734 iovss.n2560 iovss.n1450 0.00818093
R13735 iovss.n2457 iovss.n2456 0.00818093
R13736 iovss.n2449 iovss.n2448 0.00818093
R13737 iovss.n2441 iovss.n2440 0.00818093
R13738 iovss.n2473 iovss.n2472 0.00818093
R13739 iovss.n2481 iovss.n2480 0.00818093
R13740 iovss.n2424 iovss.n2423 0.00818093
R13741 iovss.n2416 iovss.n2415 0.00818093
R13742 iovss.n2497 iovss.n2496 0.00818093
R13743 iovss.n2505 iovss.n2504 0.00818093
R13744 iovss.n2456 iovss.n2455 0.00818093
R13745 iovss.n2460 iovss.n2459 0.00818093
R13746 iovss.n2450 iovss.n2449 0.00818093
R13747 iovss.n2446 iovss.n2445 0.00818093
R13748 iovss.n2442 iovss.n2441 0.00818093
R13749 iovss.n2438 iovss.n2427 0.00818093
R13750 iovss.n2472 iovss.n2471 0.00818093
R13751 iovss.n2476 iovss.n2475 0.00818093
R13752 iovss.n2480 iovss.n2479 0.00818093
R13753 iovss.n2484 iovss.n2483 0.00818093
R13754 iovss.n2425 iovss.n2424 0.00818093
R13755 iovss.n2421 iovss.n2420 0.00818093
R13756 iovss.n2417 iovss.n2416 0.00818093
R13757 iovss.n2413 iovss.n2403 0.00818093
R13758 iovss.n2496 iovss.n2495 0.00818093
R13759 iovss.n2500 iovss.n2499 0.00818093
R13760 iovss.n2506 iovss.n2505 0.00818093
R13761 iovss.n2510 iovss.n2509 0.00818093
R13762 iovss.n2040 iovss.n2039 0.00783333
R13763 iovss.n2046 iovss.n2040 0.00783333
R13764 iovss.n2047 iovss.n2046 0.00783333
R13765 iovss.n2048 iovss.n2047 0.00783333
R13766 iovss.n2049 iovss.n2048 0.00783333
R13767 iovss.n2051 iovss.n2049 0.00783333
R13768 iovss.n2051 iovss.n2050 0.00783333
R13769 iovss.n2050 iovss.n1509 0.00783333
R13770 iovss.n1510 iovss.n1509 0.00783333
R13771 iovss.n1511 iovss.n1510 0.00783333
R13772 iovss.n1517 iovss.n1511 0.00783333
R13773 iovss.n1518 iovss.n1517 0.00783333
R13774 iovss.n1519 iovss.n1518 0.00783333
R13775 iovss.n1520 iovss.n1519 0.00783333
R13776 iovss.n1525 iovss.n1520 0.00783333
R13777 iovss.n1526 iovss.n1525 0.00783333
R13778 iovss.n1527 iovss.n1526 0.00783333
R13779 iovss.n1528 iovss.n1527 0.00783333
R13780 iovss.n2406 iovss.n1528 0.00783333
R13781 iovss.n2407 iovss.n2406 0.00783333
R13782 iovss.n2408 iovss.n2407 0.00783333
R13783 iovss.n2409 iovss.n2408 0.00783333
R13784 iovss.n2430 iovss.n2409 0.00783333
R13785 iovss.n2431 iovss.n2430 0.00783333
R13786 iovss.n2432 iovss.n2431 0.00783333
R13787 iovss.n2433 iovss.n2432 0.00783333
R13788 iovss.n2434 iovss.n2433 0.00783333
R13789 iovss.n2434 iovss.n1430 0.00783333
R13790 iovss.n2591 iovss.n1430 0.00783333
R13791 iovss.n2592 iovss.n2591 0.00783333
R13792 iovss.n1504 iovss.n1484 0.00783333
R13793 iovss.n2420 iovss.n2419 0.00783333
R13794 iovss.n1504 iovss.n1451 0.00754
R13795 iovss.n2419 iovss.n2418 0.00754
R13796 iovss.n3133 iovss.n927 0.00748413
R13797 iovss.n3077 iovss.n3075 0.00748413
R13798 iovss.n3133 iovss.n3132 0.00748413
R13799 iovss.n3107 iovss.n1107 0.00748413
R13800 iovss.n2213 iovss.n2163 0.00740196
R13801 iovss.n2213 iovss.n2212 0.00740196
R13802 iovss.n2212 iovss.n2210 0.00740196
R13803 iovss.n2210 iovss.n2208 0.00740196
R13804 iovss.n2208 iovss.n2206 0.00740196
R13805 iovss.n2206 iovss.n2204 0.00740196
R13806 iovss.n2204 iovss.n2202 0.00740196
R13807 iovss.n2202 iovss.n1890 0.00740196
R13808 iovss.n2245 iovss.n1890 0.00740196
R13809 iovss.n2245 iovss.n1872 0.00740196
R13810 iovss.n2287 iovss.n1872 0.00740196
R13811 iovss.n2287 iovss.n2286 0.00740196
R13812 iovss.n2286 iovss.n2284 0.00740196
R13813 iovss.n2284 iovss.n2282 0.00740196
R13814 iovss.n2282 iovss.n2280 0.00740196
R13815 iovss.n2280 iovss.n2278 0.00740196
R13816 iovss.n2278 iovss.n2276 0.00740196
R13817 iovss.n2276 iovss.n2274 0.00740196
R13818 iovss.n2274 iovss.n1703 0.00740196
R13819 iovss.n2294 iovss.n1703 0.00740196
R13820 iovss.n2295 iovss.n2294 0.00740196
R13821 iovss.n2297 iovss.n2295 0.00740196
R13822 iovss.n2297 iovss.n1696 0.00740196
R13823 iovss.n2308 iovss.n1696 0.00740196
R13824 iovss.n2310 iovss.n2308 0.00740196
R13825 iovss.n2312 iovss.n2310 0.00740196
R13826 iovss.n2312 iovss.n1688 0.00740196
R13827 iovss.n2326 iovss.n1688 0.00740196
R13828 iovss.n2328 iovss.n2326 0.00740196
R13829 iovss.n2328 iovss.n1678 0.00740196
R13830 iovss.n2353 iovss.n1678 0.00740196
R13831 iovss.n2353 iovss.n2352 0.00740196
R13832 iovss.n2352 iovss.n2351 0.00740196
R13833 iovss.n2351 iovss.n1220 0.00740196
R13834 iovss.n3082 iovss.n1220 0.00740196
R13835 iovss.n3082 iovss.n3081 0.00740196
R13836 iovss.n3081 iovss.n1223 0.00740196
R13837 iovss.n2293 iovss.n1652 0.00740196
R13838 iovss.n2354 iovss.n1677 0.00740196
R13839 iovss.n276 iovss.n254 0.00740196
R13840 iovss.n945 iovss.n867 0.00740196
R13841 iovss.n3244 iovss.n769 0.00740196
R13842 iovss.n3244 iovss.n771 0.00740196
R13843 iovss.n3237 iovss.n771 0.00740196
R13844 iovss.n3237 iovss.n3236 0.00740196
R13845 iovss.n3236 iovss.n784 0.00740196
R13846 iovss.n3229 iovss.n784 0.00740196
R13847 iovss.n3229 iovss.n3228 0.00740196
R13848 iovss.n3228 iovss.n794 0.00740196
R13849 iovss.n3221 iovss.n794 0.00740196
R13850 iovss.n3221 iovss.n3220 0.00740196
R13851 iovss.n3220 iovss.n802 0.00740196
R13852 iovss.n3213 iovss.n802 0.00740196
R13853 iovss.n3213 iovss.n3212 0.00740196
R13854 iovss.n3212 iovss.n812 0.00740196
R13855 iovss.n3205 iovss.n812 0.00740196
R13856 iovss.n3205 iovss.n3204 0.00740196
R13857 iovss.n3204 iovss.n822 0.00740196
R13858 iovss.n3197 iovss.n822 0.00740196
R13859 iovss.n3197 iovss.n3196 0.00740196
R13860 iovss.n3196 iovss.n831 0.00740196
R13861 iovss.n3189 iovss.n831 0.00740196
R13862 iovss.n3189 iovss.n3188 0.00740196
R13863 iovss.n3188 iovss.n840 0.00740196
R13864 iovss.n3181 iovss.n840 0.00740196
R13865 iovss.n3181 iovss.n3180 0.00740196
R13866 iovss.n3180 iovss.n849 0.00740196
R13867 iovss.n3173 iovss.n849 0.00740196
R13868 iovss.n3173 iovss.n3172 0.00740196
R13869 iovss.n3172 iovss.n859 0.00740196
R13870 iovss.n3165 iovss.n859 0.00740196
R13871 iovss.n3165 iovss.n3164 0.00740196
R13872 iovss.n3164 iovss.n868 0.00740196
R13873 iovss.n3157 iovss.n868 0.00740196
R13874 iovss.n3157 iovss.n3156 0.00740196
R13875 iovss.n3156 iovss.n877 0.00740196
R13876 iovss.n3149 iovss.n877 0.00740196
R13877 iovss.n3149 iovss.n3148 0.00740196
R13878 iovss.n1111 iovss 0.00727871
R13879 iovss.n3107 iovss.n3106 0.00727735
R13880 iovss.n3462 iovss 0.0071
R13881 iovss.n2072 iovss.n2038 0.00694773
R13882 iovss.n2594 iovss.n2593 0.00694773
R13883 iovss.n2929 iovss 0.00671176
R13884 iovss.n2930 iovss.n904 0.00666247
R13885 iovss.n2562 iovss.n2540 0.00666
R13886 iovss.n2485 iovss.n2484 0.00666
R13887 iovss.n1416 iovss 0.00666
R13888 iovss.n2355 iovss.n2354 0.00653922
R13889 iovss.n867 iovss.n219 0.00653922
R13890 iovss.n2532 iovss.n1453 0.00636667
R13891 iovss.n2494 iovss.n2493 0.00636667
R13892 iovss.n3077 iovss.n904 0.00627731
R13893 iovss.n2290 iovss.n1871 0.00619412
R13894 iovss.n3392 iovss.n332 0.00619412
R13895 iovss.n2078 iovss.n2077 0.00607333
R13896 iovss.n1425 iovss.n1415 0.00607333
R13897 iovss.n595 iovss.n552 0.00578
R13898 iovss.n1057 iovss.n904 0.0057381
R13899 iovss.n2931 iovss.n904 0.0057381
R13900 iovss.n3277 iovss.n423 0.00567
R13901 iovss.n473 iovss.n419 0.00567
R13902 iovss.n1137 iovss.n904 0.00565631
R13903 iovss.n593 iovss.n547 0.00556
R13904 iovss.n1996 iovss.n1985 0.00548667
R13905 iovss.n2477 iovss.n2476 0.00548667
R13906 iovss.n3328 iovss.n126 0.00545
R13907 iovss.n3325 iovss.n135 0.00545
R13908 iovss.n558 iovss.n555 0.00534
R13909 iovss.n3275 iovss.n425 0.00523
R13910 iovss.n3288 iovss.n417 0.00523
R13911 iovss.n2530 iovss.n1455 0.00519333
R13912 iovss.n2503 iovss.n2501 0.00519333
R13913 iovss.n567 iovss.n544 0.00512
R13914 iovss.n3330 iovss.n122 0.00501
R13915 iovss.n3323 iovss.n138 0.00501
R13916 iovss.n586 iovss.n572 0.005
R13917 iovss.n586 iovss.n570 0.005
R13918 iovss.n590 iovss.n570 0.005
R13919 iovss.n590 iovss.n565 0.005
R13920 iovss.n600 iovss.n565 0.005
R13921 iovss.n600 iovss.n563 0.005
R13922 iovss.n604 iovss.n563 0.005
R13923 iovss.n604 iovss.n485 0.005
R13924 iovss.n3265 iovss.n485 0.005
R13925 iovss.n3265 iovss.n483 0.005
R13926 iovss.n3269 iovss.n483 0.005
R13927 iovss.n3269 iovss.n478 0.005
R13928 iovss.n3281 iovss.n478 0.005
R13929 iovss.n3281 iovss.n476 0.005
R13930 iovss.n3285 iovss.n476 0.005
R13931 iovss.n3285 iovss.n471 0.005
R13932 iovss.n3296 iovss.n471 0.005
R13933 iovss.n3296 iovss.n469 0.005
R13934 iovss.n3301 iovss.n469 0.005
R13935 iovss.n3303 iovss.n3301 0.005
R13936 iovss.n3305 iovss.n3303 0.005
R13937 iovss.n3305 iovss.n467 0.005
R13938 iovss.n3310 iovss.n467 0.005
R13939 iovss.n3312 iovss.n3310 0.005
R13940 iovss.n3314 iovss.n3312 0.005
R13941 iovss.n3314 iovss.n464 0.005
R13942 iovss.n3318 iovss.n464 0.005
R13943 iovss.n3318 iovss.n75 0.005
R13944 iovss.n3442 iovss.n75 0.005
R13945 iovss.n3442 iovss.n72 0.005
R13946 iovss.n3447 iovss.n72 0.005
R13947 iovss.n3447 iovss.n73 0.005
R13948 iovss.n73 iovss.n65 0.005
R13949 iovss.n3459 iovss.n65 0.005
R13950 iovss.n3459 iovss.n63 0.005
R13951 iovss.n3463 iovss.n63 0.005
R13952 iovss.n2074 iovss.n2032 0.0049
R13953 iovss.n2598 iovss.n2597 0.0049
R13954 iovss.n588 iovss.n587 0.0049
R13955 iovss.n589 iovss.n588 0.0049
R13956 iovss.n589 iovss.n564 0.0049
R13957 iovss.n601 iovss.n564 0.0049
R13958 iovss.n602 iovss.n601 0.0049
R13959 iovss.n603 iovss.n602 0.0049
R13960 iovss.n603 iovss.n484 0.0049
R13961 iovss.n3266 iovss.n484 0.0049
R13962 iovss.n3267 iovss.n3266 0.0049
R13963 iovss.n3268 iovss.n3267 0.0049
R13964 iovss.n3268 iovss.n477 0.0049
R13965 iovss.n3282 iovss.n477 0.0049
R13966 iovss.n3283 iovss.n3282 0.0049
R13967 iovss.n3284 iovss.n3283 0.0049
R13968 iovss.n3284 iovss.n470 0.0049
R13969 iovss.n3297 iovss.n470 0.0049
R13970 iovss.n3298 iovss.n3297 0.0049
R13971 iovss.n3299 iovss.n3298 0.0049
R13972 iovss.n3299 iovss.n468 0.0049
R13973 iovss.n3306 iovss.n468 0.0049
R13974 iovss.n3307 iovss.n3306 0.0049
R13975 iovss.n3308 iovss.n3307 0.0049
R13976 iovss.n3308 iovss.n465 0.0049
R13977 iovss.n3315 iovss.n465 0.0049
R13978 iovss.n3316 iovss.n3315 0.0049
R13979 iovss.n3317 iovss.n3316 0.0049
R13980 iovss.n3317 iovss.n74 0.0049
R13981 iovss.n3443 iovss.n74 0.0049
R13982 iovss.n3444 iovss.n3443 0.0049
R13983 iovss.n3446 iovss.n3444 0.0049
R13984 iovss.n3446 iovss.n3445 0.0049
R13985 iovss.n3445 iovss.n64 0.0049
R13986 iovss.n3460 iovss.n64 0.0049
R13987 iovss.n3461 iovss.n3460 0.0049
R13988 iovss.n3462 iovss.n3461 0.0049
R13989 iovss.n609 iovss.n608 0.0049
R13990 iovss.n26 iovss.n1 0.00479417
R13991 iovss.n43 iovss.n2 0.00479417
R13992 iovss.n27 iovss.n2 0.00479417
R13993 iovss.n34 iovss.n13 0.00479417
R13994 iovss.n42 iovss.n12 0.00479417
R13995 iovss.n33 iovss.n12 0.00479417
R13996 iovss.n28 iovss.n4 0.00479417
R13997 iovss.n41 iovss.n5 0.00479417
R13998 iovss.n29 iovss.n5 0.00479417
R13999 iovss.n32 iovss.n6 0.00479417
R14000 iovss.n40 iovss.n9 0.00479417
R14001 iovss.n30 iovss.n7 0.00479417
R14002 iovss.n39 iovss.n8 0.00479417
R14003 iovss.n3476 iovss.n3471 0.00479417
R14004 iovss.n3479 iovss.n15 0.00479417
R14005 iovss.n3476 iovss.n15 0.00479417
R14006 iovss.n3471 iovss.n8 0.00479417
R14007 iovss.n39 iovss.n7 0.00479417
R14008 iovss.n30 iovss.n9 0.00479417
R14009 iovss.n32 iovss.n10 0.00479417
R14010 iovss.n29 iovss.n10 0.00479417
R14011 iovss.n41 iovss.n11 0.00479417
R14012 iovss.n28 iovss.n11 0.00479417
R14013 iovss.n33 iovss.n4 0.00479417
R14014 iovss.n42 iovss.n3 0.00479417
R14015 iovss.n34 iovss.n3 0.00479417
R14016 iovss.n27 iovss.n13 0.00479417
R14017 iovss.n43 iovss.n14 0.00479417
R14018 iovss.n26 iovss.n14 0.00479417
R14019 iovss.n40 iovss.n6 0.00479417
R14020 iovss.n3273 iovss.n427 0.00479
R14021 iovss.n3290 iovss.n415 0.00479
R14022 iovss.n3080 iovss.n3079 0.0047102
R14023 iovss.n3144 iovss.n885 0.0047102
R14024 iovss.n582 iovss.n541 0.00468
R14025 iovss.n3321 iovss.n141 0.00457
R14026 iovss.n613 iovss.n612 0.00446
R14027 iovss.n2163 iovss.n2161 0.00442211
R14028 iovss.n769 iovss.n732 0.00442211
R14029 iovss iovss.n3480 0.004405
R14030 iovss.n3343 iovss.n388 0.00435
R14031 iovss.n452 iovss.n413 0.00435
R14032 iovss.n2054 iovss.n2017 0.00431333
R14033 iovss.n2469 iovss.n2427 0.00431333
R14034 iovss.n580 iovss.n538 0.00424
R14035 iovss.n145 iovss.n144 0.00413
R14036 iovss.n2528 iovss.n1457 0.00402
R14037 iovss.n2511 iovss.n1547 0.00402
R14038 iovss.n3260 iovss.n3259 0.00402
R14039 iovss.n3465 iovss.n17 0.003965
R14040 iovss.n2178 iovss.n2177 0.00395098
R14041 iovss.n2179 iovss.n2178 0.00395098
R14042 iovss.n2179 iovss.n2164 0.00395098
R14043 iovss.n2181 iovss.n2164 0.00395098
R14044 iovss.n2181 iovss.n2165 0.00395098
R14045 iovss.n2174 iovss.n2165 0.00395098
R14046 iovss.n2174 iovss.n2166 0.00395098
R14047 iovss.n2186 iovss.n2166 0.00395098
R14048 iovss.n2186 iovss.n2167 0.00395098
R14049 iovss.n2188 iovss.n2167 0.00395098
R14050 iovss.n2188 iovss.n2168 0.00395098
R14051 iovss.n2190 iovss.n2168 0.00395098
R14052 iovss.n2190 iovss.n2169 0.00395098
R14053 iovss.n2170 iovss.n2169 0.00395098
R14054 iovss.n2200 iovss.n2170 0.00395098
R14055 iovss.n2200 iovss.n2199 0.00395098
R14056 iovss.n2199 iovss.n2171 0.00395098
R14057 iovss.n2171 iovss.n1889 0.00395098
R14058 iovss.n2246 iovss.n1889 0.00395098
R14059 iovss.n2247 iovss.n2246 0.00395098
R14060 iovss.n2248 iovss.n2247 0.00395098
R14061 iovss.n2249 iovss.n2248 0.00395098
R14062 iovss.n2249 iovss.n1873 0.00395098
R14063 iovss.n2251 iovss.n1873 0.00395098
R14064 iovss.n2251 iovss.n1874 0.00395098
R14065 iovss.n2253 iovss.n1874 0.00395098
R14066 iovss.n2253 iovss.n1875 0.00395098
R14067 iovss.n1884 iovss.n1875 0.00395098
R14068 iovss.n1884 iovss.n1876 0.00395098
R14069 iovss.n2258 iovss.n1876 0.00395098
R14070 iovss.n2258 iovss.n1877 0.00395098
R14071 iovss.n2260 iovss.n1877 0.00395098
R14072 iovss.n2260 iovss.n1878 0.00395098
R14073 iovss.n2262 iovss.n1878 0.00395098
R14074 iovss.n2262 iovss.n1879 0.00395098
R14075 iovss.n1880 iovss.n1879 0.00395098
R14076 iovss.n2272 iovss.n1880 0.00395098
R14077 iovss.n2272 iovss.n2271 0.00395098
R14078 iovss.n2271 iovss.n1881 0.00395098
R14079 iovss.n2268 iovss.n1881 0.00395098
R14080 iovss.n2268 iovss.n1705 0.00395098
R14081 iovss.n1705 iovss.n1704 0.00395098
R14082 iovss.n1704 iovss.n1701 0.00395098
R14083 iovss.n2299 iovss.n1701 0.00395098
R14084 iovss.n2299 iovss.n2298 0.00395098
R14085 iovss.n2298 iovss.n1702 0.00395098
R14086 iovss.n1702 iovss.n1697 0.00395098
R14087 iovss.n2305 iovss.n1697 0.00395098
R14088 iovss.n2307 iovss.n2305 0.00395098
R14089 iovss.n2307 iovss.n2306 0.00395098
R14090 iovss.n2306 iovss.n1693 0.00395098
R14091 iovss.n2314 iovss.n1693 0.00395098
R14092 iovss.n2314 iovss.n2313 0.00395098
R14093 iovss.n2313 iovss.n1694 0.00395098
R14094 iovss.n1694 iovss.n1689 0.00395098
R14095 iovss.n2323 iovss.n1689 0.00395098
R14096 iovss.n2324 iovss.n2323 0.00395098
R14097 iovss.n2324 iovss.n1686 0.00395098
R14098 iovss.n2329 iovss.n1686 0.00395098
R14099 iovss.n2330 iovss.n2329 0.00395098
R14100 iovss.n2331 iovss.n2330 0.00395098
R14101 iovss.n2332 iovss.n2331 0.00395098
R14102 iovss.n2332 iovss.n1679 0.00395098
R14103 iovss.n2334 iovss.n1679 0.00395098
R14104 iovss.n2334 iovss.n1680 0.00395098
R14105 iovss.n1681 iovss.n1680 0.00395098
R14106 iovss.n2350 iovss.n1681 0.00395098
R14107 iovss.n2350 iovss.n2349 0.00395098
R14108 iovss.n2349 iovss.n1682 0.00395098
R14109 iovss.n2346 iovss.n1682 0.00395098
R14110 iovss.n2346 iovss.n1221 0.00395098
R14111 iovss.n2344 iovss.n1221 0.00395098
R14112 iovss.n2344 iovss.n1222 0.00395098
R14113 iovss.n2342 iovss.n1222 0.00395098
R14114 iovss.n776 iovss.n775 0.00395098
R14115 iovss.n775 iovss.n772 0.00395098
R14116 iovss.n3243 iovss.n772 0.00395098
R14117 iovss.n3243 iovss.n3242 0.00395098
R14118 iovss.n3242 iovss.n773 0.00395098
R14119 iovss.n3239 iovss.n773 0.00395098
R14120 iovss.n3239 iovss.n3238 0.00395098
R14121 iovss.n3238 iovss.n781 0.00395098
R14122 iovss.n3235 iovss.n781 0.00395098
R14123 iovss.n3235 iovss.n3234 0.00395098
R14124 iovss.n3234 iovss.n785 0.00395098
R14125 iovss.n3231 iovss.n785 0.00395098
R14126 iovss.n3231 iovss.n3230 0.00395098
R14127 iovss.n3230 iovss.n790 0.00395098
R14128 iovss.n3227 iovss.n790 0.00395098
R14129 iovss.n3227 iovss.n3226 0.00395098
R14130 iovss.n3226 iovss.n795 0.00395098
R14131 iovss.n3223 iovss.n795 0.00395098
R14132 iovss.n3223 iovss.n3222 0.00395098
R14133 iovss.n3222 iovss.n800 0.00395098
R14134 iovss.n3219 iovss.n800 0.00395098
R14135 iovss.n3219 iovss.n3218 0.00395098
R14136 iovss.n3218 iovss.n803 0.00395098
R14137 iovss.n3215 iovss.n803 0.00395098
R14138 iovss.n3215 iovss.n3214 0.00395098
R14139 iovss.n3214 iovss.n808 0.00395098
R14140 iovss.n3211 iovss.n808 0.00395098
R14141 iovss.n3211 iovss.n3210 0.00395098
R14142 iovss.n3210 iovss.n813 0.00395098
R14143 iovss.n3207 iovss.n813 0.00395098
R14144 iovss.n3207 iovss.n3206 0.00395098
R14145 iovss.n3206 iovss.n818 0.00395098
R14146 iovss.n3203 iovss.n818 0.00395098
R14147 iovss.n3203 iovss.n3202 0.00395098
R14148 iovss.n3202 iovss.n823 0.00395098
R14149 iovss.n3199 iovss.n823 0.00395098
R14150 iovss.n3199 iovss.n3198 0.00395098
R14151 iovss.n3198 iovss.n828 0.00395098
R14152 iovss.n3195 iovss.n828 0.00395098
R14153 iovss.n3195 iovss.n3194 0.00395098
R14154 iovss.n3194 iovss.n832 0.00395098
R14155 iovss.n3191 iovss.n832 0.00395098
R14156 iovss.n3191 iovss.n3190 0.00395098
R14157 iovss.n3190 iovss.n837 0.00395098
R14158 iovss.n3187 iovss.n837 0.00395098
R14159 iovss.n3187 iovss.n3186 0.00395098
R14160 iovss.n3186 iovss.n841 0.00395098
R14161 iovss.n3183 iovss.n841 0.00395098
R14162 iovss.n3183 iovss.n3182 0.00395098
R14163 iovss.n3182 iovss.n846 0.00395098
R14164 iovss.n3179 iovss.n846 0.00395098
R14165 iovss.n3179 iovss.n3178 0.00395098
R14166 iovss.n3178 iovss.n850 0.00395098
R14167 iovss.n3175 iovss.n850 0.00395098
R14168 iovss.n3175 iovss.n3174 0.00395098
R14169 iovss.n3174 iovss.n855 0.00395098
R14170 iovss.n3171 iovss.n855 0.00395098
R14171 iovss.n3171 iovss.n3170 0.00395098
R14172 iovss.n3170 iovss.n860 0.00395098
R14173 iovss.n3167 iovss.n860 0.00395098
R14174 iovss.n3167 iovss.n3166 0.00395098
R14175 iovss.n3166 iovss.n865 0.00395098
R14176 iovss.n3163 iovss.n865 0.00395098
R14177 iovss.n3163 iovss.n3162 0.00395098
R14178 iovss.n3162 iovss.n869 0.00395098
R14179 iovss.n3159 iovss.n869 0.00395098
R14180 iovss.n3159 iovss.n3158 0.00395098
R14181 iovss.n3158 iovss.n874 0.00395098
R14182 iovss.n3155 iovss.n874 0.00395098
R14183 iovss.n3155 iovss.n3154 0.00395098
R14184 iovss.n3154 iovss.n878 0.00395098
R14185 iovss.n3151 iovss.n878 0.00395098
R14186 iovss.n3151 iovss.n3150 0.00395098
R14187 iovss.n3150 iovss.n884 0.00395098
R14188 iovss.n3338 iovss.n362 0.00391
R14189 iovss.n3083 iovss.n1219 0.00384745
R14190 iovss.n2773 iovss.n914 0.00384745
R14191 iovss.n2035 iovss.n2030 0.00372667
R14192 iovss.n2581 iovss.n2580 0.00372667
R14193 iovss.n631 iovss.n538 0.00369419
R14194 iovss.n630 iovss.n540 0.00369419
R14195 iovss.n539 iovss.n535 0.00369419
R14196 iovss.n629 iovss.n541 0.00369419
R14197 iovss.n628 iovss.n543 0.00369419
R14198 iovss.n542 iovss.n533 0.00369419
R14199 iovss.n627 iovss.n544 0.00369419
R14200 iovss.n626 iovss.n546 0.00369419
R14201 iovss.n545 iovss.n531 0.00369419
R14202 iovss.n625 iovss.n547 0.00369419
R14203 iovss.n548 iovss.n530 0.00369419
R14204 iovss.n624 iovss.n529 0.00369419
R14205 iovss.n550 iovss.n529 0.00369419
R14206 iovss.n623 iovss.n528 0.00369419
R14207 iovss.n622 iovss.n527 0.00369419
R14208 iovss.n553 iovss.n527 0.00369419
R14209 iovss.n621 iovss.n526 0.00369419
R14210 iovss.n620 iovss.n525 0.00369419
R14211 iovss.n556 iovss.n525 0.00369419
R14212 iovss.n619 iovss.n524 0.00369419
R14213 iovss.n618 iovss.n523 0.00369419
R14214 iovss.n610 iovss.n523 0.00369419
R14215 iovss.n617 iovss.n522 0.00369419
R14216 iovss.n616 iovss.n521 0.00369419
R14217 iovss.n3256 iovss.n521 0.00369419
R14218 iovss.n3255 iovss.n489 0.00369419
R14219 iovss.n518 iovss.n497 0.00369419
R14220 iovss.n519 iovss.n518 0.00369419
R14221 iovss.n428 iovss.n379 0.00369419
R14222 iovss.n430 iovss.n428 0.00369419
R14223 iovss.n427 iovss.n378 0.00369419
R14224 iovss.n426 iovss.n377 0.00369419
R14225 iovss.n433 iovss.n426 0.00369419
R14226 iovss.n425 iovss.n376 0.00369419
R14227 iovss.n424 iovss.n375 0.00369419
R14228 iovss.n436 iovss.n424 0.00369419
R14229 iovss.n423 iovss.n374 0.00369419
R14230 iovss.n422 iovss.n421 0.00369419
R14231 iovss.n439 iovss.n372 0.00369419
R14232 iovss.n438 iovss.n420 0.00369419
R14233 iovss.n440 iovss.n371 0.00369419
R14234 iovss.n442 iovss.n370 0.00369419
R14235 iovss.n441 iovss.n418 0.00369419
R14236 iovss.n443 iovss.n369 0.00369419
R14237 iovss.n445 iovss.n368 0.00369419
R14238 iovss.n444 iovss.n416 0.00369419
R14239 iovss.n446 iovss.n367 0.00369419
R14240 iovss.n448 iovss.n366 0.00369419
R14241 iovss.n447 iovss.n414 0.00369419
R14242 iovss.n449 iovss.n365 0.00369419
R14243 iovss.n451 iovss.n364 0.00369419
R14244 iovss.n450 iovss.n412 0.00369419
R14245 iovss.n3339 iovss.n363 0.00369419
R14246 iovss.n3340 iovss.n362 0.00369419
R14247 iovss.n409 iovss.n361 0.00369419
R14248 iovss.n410 iovss.n409 0.00369419
R14249 iovss.n170 iovss.n120 0.00369419
R14250 iovss.n163 iovss.n118 0.00369419
R14251 iovss.n121 iovss.n118 0.00369419
R14252 iovss.n123 iovss.n117 0.00369419
R14253 iovss.n162 iovss.n116 0.00369419
R14254 iovss.n125 iovss.n116 0.00369419
R14255 iovss.n127 iovss.n115 0.00369419
R14256 iovss.n161 iovss.n114 0.00369419
R14257 iovss.n129 iovss.n114 0.00369419
R14258 iovss.n160 iovss.n113 0.00369419
R14259 iovss.n131 iovss.n113 0.00369419
R14260 iovss.n159 iovss.n112 0.00369419
R14261 iovss.n133 iovss.n112 0.00369419
R14262 iovss.n158 iovss.n111 0.00369419
R14263 iovss.n157 iovss.n110 0.00369419
R14264 iovss.n136 iovss.n110 0.00369419
R14265 iovss.n156 iovss.n109 0.00369419
R14266 iovss.n155 iovss.n108 0.00369419
R14267 iovss.n139 iovss.n108 0.00369419
R14268 iovss.n154 iovss.n107 0.00369419
R14269 iovss.n153 iovss.n106 0.00369419
R14270 iovss.n142 iovss.n106 0.00369419
R14271 iovss.n152 iovss.n105 0.00369419
R14272 iovss.n151 iovss.n104 0.00369419
R14273 iovss.n146 iovss.n104 0.00369419
R14274 iovss.n150 iovss.n78 0.00369419
R14275 iovss.n103 iovss.n86 0.00369419
R14276 iovss.n3433 iovss.n103 0.00369419
R14277 iovss.n148 iovss.n101 0.00369419
R14278 iovss.n3477 iovss.n20 0.00369419
R14279 iovss.n51 iovss.n50 0.00369419
R14280 iovss.n3475 iovss.n19 0.00369419
R14281 iovss.n3474 iovss.n18 0.00369419
R14282 iovss.n54 iovss.n53 0.00369419
R14283 iovss.n3473 iovss.n17 0.00369419
R14284 iovss.n3472 iovss.n16 0.00369419
R14285 iovss.n57 iovss.n56 0.00369419
R14286 iovss.n3480 iovss.n0 0.00369419
R14287 iovss.n631 iovss.n537 0.00369419
R14288 iovss.n630 iovss.n536 0.00369419
R14289 iovss.n629 iovss.n535 0.00369419
R14290 iovss.n628 iovss.n534 0.00369419
R14291 iovss.n627 iovss.n533 0.00369419
R14292 iovss.n626 iovss.n532 0.00369419
R14293 iovss.n625 iovss.n531 0.00369419
R14294 iovss.n624 iovss.n549 0.00369419
R14295 iovss.n623 iovss.n551 0.00369419
R14296 iovss.n622 iovss.n552 0.00369419
R14297 iovss.n621 iovss.n554 0.00369419
R14298 iovss.n620 iovss.n555 0.00369419
R14299 iovss.n619 iovss.n557 0.00369419
R14300 iovss.n618 iovss.n609 0.00369419
R14301 iovss.n617 iovss.n611 0.00369419
R14302 iovss.n616 iovss.n613 0.00369419
R14303 iovss.n3257 iovss.n3255 0.00369419
R14304 iovss.n3259 iovss.n497 0.00369419
R14305 iovss.n540 iovss.n539 0.00369419
R14306 iovss.n543 iovss.n542 0.00369419
R14307 iovss.n546 iovss.n545 0.00369419
R14308 iovss.n549 iovss.n548 0.00369419
R14309 iovss.n551 iovss.n550 0.00369419
R14310 iovss.n554 iovss.n553 0.00369419
R14311 iovss.n557 iovss.n556 0.00369419
R14312 iovss.n611 iovss.n610 0.00369419
R14313 iovss.n3257 iovss.n3256 0.00369419
R14314 iovss.n614 iovss.n519 0.00369419
R14315 iovss.n429 iovss.n379 0.00369419
R14316 iovss.n431 iovss.n378 0.00369419
R14317 iovss.n432 iovss.n377 0.00369419
R14318 iovss.n434 iovss.n376 0.00369419
R14319 iovss.n435 iovss.n375 0.00369419
R14320 iovss.n437 iovss.n374 0.00369419
R14321 iovss.n422 iovss.n372 0.00369419
R14322 iovss.n420 iovss.n371 0.00369419
R14323 iovss.n419 iovss.n370 0.00369419
R14324 iovss.n418 iovss.n369 0.00369419
R14325 iovss.n417 iovss.n368 0.00369419
R14326 iovss.n416 iovss.n367 0.00369419
R14327 iovss.n415 iovss.n366 0.00369419
R14328 iovss.n414 iovss.n365 0.00369419
R14329 iovss.n413 iovss.n364 0.00369419
R14330 iovss.n412 iovss.n363 0.00369419
R14331 iovss.n3341 iovss.n361 0.00369419
R14332 iovss.n431 iovss.n430 0.00369419
R14333 iovss.n434 iovss.n433 0.00369419
R14334 iovss.n437 iovss.n436 0.00369419
R14335 iovss.n421 iovss.n373 0.00369419
R14336 iovss.n439 iovss.n438 0.00369419
R14337 iovss.n442 iovss.n441 0.00369419
R14338 iovss.n445 iovss.n444 0.00369419
R14339 iovss.n448 iovss.n447 0.00369419
R14340 iovss.n451 iovss.n450 0.00369419
R14341 iovss.n3341 iovss.n3340 0.00369419
R14342 iovss.n3333 iovss.n410 0.00369419
R14343 iovss.n3478 iovss.n3477 0.00369419
R14344 iovss.n3475 iovss.n51 0.00369419
R14345 iovss.n3474 iovss.n52 0.00369419
R14346 iovss.n3473 iovss.n54 0.00369419
R14347 iovss.n3472 iovss.n55 0.00369419
R14348 iovss.n57 iovss.n0 0.00369419
R14349 iovss.n50 iovss.n20 0.00369419
R14350 iovss.n53 iovss.n18 0.00369419
R14351 iovss.n56 iovss.n16 0.00369419
R14352 iovss.n163 iovss.n120 0.00369419
R14353 iovss.n162 iovss.n124 0.00369419
R14354 iovss.n161 iovss.n128 0.00369419
R14355 iovss.n160 iovss.n130 0.00369419
R14356 iovss.n159 iovss.n132 0.00369419
R14357 iovss.n158 iovss.n134 0.00369419
R14358 iovss.n157 iovss.n135 0.00369419
R14359 iovss.n156 iovss.n137 0.00369419
R14360 iovss.n155 iovss.n138 0.00369419
R14361 iovss.n154 iovss.n140 0.00369419
R14362 iovss.n153 iovss.n141 0.00369419
R14363 iovss.n152 iovss.n143 0.00369419
R14364 iovss.n151 iovss.n145 0.00369419
R14365 iovss.n150 iovss.n147 0.00369419
R14366 iovss.n3436 iovss.n86 0.00369419
R14367 iovss.n171 iovss.n170 0.00369419
R14368 iovss.n122 iovss.n121 0.00369419
R14369 iovss.n124 iovss.n123 0.00369419
R14370 iovss.n126 iovss.n125 0.00369419
R14371 iovss.n128 iovss.n127 0.00369419
R14372 iovss.n130 iovss.n129 0.00369419
R14373 iovss.n132 iovss.n131 0.00369419
R14374 iovss.n134 iovss.n133 0.00369419
R14375 iovss.n137 iovss.n136 0.00369419
R14376 iovss.n140 iovss.n139 0.00369419
R14377 iovss.n143 iovss.n142 0.00369419
R14378 iovss.n147 iovss.n146 0.00369419
R14379 iovss.n3434 iovss.n148 0.00369419
R14380 iovss.n3434 iovss.n3433 0.00369419
R14381 iovss.n3437 iovss.n3436 0.00369
R14382 iovss.n3104 iovss 0.00358123
R14383 iovss.n3467 iovss.n19 0.003525
R14384 iovss.n3478 iovss.n3470 0.003305
R14385 iovss.n3109 iovss.n989 0.00326078
R14386 iovss.n3130 iovss.n875 0.00326078
R14387 iovss.n94 iovss.n68 0.00325
R14388 iovss.n572 iovss.n571 0.00324093
R14389 iovss.n3102 iovss.n3101 0.00314334
R14390 iovss.n1113 iovss.n1112 0.00314333
R14391 iovss.n2056 iovss.n2019 0.00314
R14392 iovss.n2445 iovss.n2444 0.00314
R14393 iovss.n101 iovss.n94 0.00314
R14394 iovss.n2601 iovss.n1410 0.00314
R14395 iovss.n3134 iovss.n904 0.00306909
R14396 iovss.n3098 iovss.n1116 0.00298471
R14397 iovss.n907 iovss.n876 0.00298471
R14398 iovss.n3335 iovss.n3333 0.00292
R14399 iovss.n1961 iovss.n1871 0.00291569
R14400 iovss.n672 iovss.n332 0.00291569
R14401 iovss.n3467 iovss.n52 0.002865
R14402 iovss.n1514 iovss.n1459 0.00284667
R14403 iovss.n1537 iovss.n1467 0.00284667
R14404 iovss.n2565 iovss.n2564 0.00284667
R14405 iovss.n3247 iovss.n768 0.00281579
R14406 iovss.n768 iovss.n756 0.00281579
R14407 iovss.n756 iovss.n755 0.00281579
R14408 iovss.n755 iovss.n754 0.00281579
R14409 iovss.n754 iovss.n753 0.00281579
R14410 iovss.n753 iovss.n752 0.00281579
R14411 iovss.n752 iovss.n751 0.00281579
R14412 iovss.n751 iovss.n750 0.00281579
R14413 iovss.n750 iovss.n749 0.00281579
R14414 iovss.n749 iovss.n748 0.00281579
R14415 iovss.n748 iovss.n747 0.00281579
R14416 iovss.n747 iovss.n746 0.00281579
R14417 iovss.n746 iovss.n745 0.00281579
R14418 iovss.n745 iovss.n744 0.00281579
R14419 iovss.n744 iovss.n743 0.00281579
R14420 iovss.n743 iovss.n633 0.00281579
R14421 iovss.n3252 iovss.n634 0.00281579
R14422 iovss.n693 iovss.n634 0.00281579
R14423 iovss.n709 iovss.n693 0.00281579
R14424 iovss.n709 iovss.n708 0.00281579
R14425 iovss.n708 iovss.n707 0.00281579
R14426 iovss.n707 iovss.n706 0.00281579
R14427 iovss.n706 iovss.n705 0.00281579
R14428 iovss.n705 iovss.n704 0.00281579
R14429 iovss.n704 iovss.n703 0.00281579
R14430 iovss.n703 iovss.n702 0.00281579
R14431 iovss.n702 iovss.n701 0.00281579
R14432 iovss.n701 iovss.n700 0.00281579
R14433 iovss.n700 iovss.n699 0.00281579
R14434 iovss.n699 iovss.n698 0.00281579
R14435 iovss.n698 iovss.n697 0.00281579
R14436 iovss.n697 iovss.n696 0.00281579
R14437 iovss.n696 iovss.n695 0.00281579
R14438 iovss.n695 iovss.n694 0.00281579
R14439 iovss.n359 iovss.n334 0.00281579
R14440 iovss.n3389 iovss.n359 0.00281579
R14441 iovss.n3389 iovss.n3388 0.00281579
R14442 iovss.n3388 iovss.n3377 0.00281579
R14443 iovss.n3377 iovss.n3376 0.00281579
R14444 iovss.n3376 iovss.n3375 0.00281579
R14445 iovss.n3375 iovss.n3374 0.00281579
R14446 iovss.n3374 iovss.n3373 0.00281579
R14447 iovss.n3373 iovss.n3372 0.00281579
R14448 iovss.n3372 iovss.n3371 0.00281579
R14449 iovss.n3371 iovss.n3370 0.00281579
R14450 iovss.n3370 iovss.n3369 0.00281579
R14451 iovss.n3369 iovss.n3368 0.00281579
R14452 iovss.n3368 iovss.n3367 0.00281579
R14453 iovss.n3367 iovss.n3366 0.00281579
R14454 iovss.n3366 iovss.n3365 0.00281579
R14455 iovss.n3365 iovss.n3364 0.00281579
R14456 iovss.n3364 iovss.n3363 0.00281579
R14457 iovss.n3361 iovss.n3360 0.00281579
R14458 iovss.n3360 iovss.n3359 0.00281579
R14459 iovss.n3359 iovss.n3358 0.00281579
R14460 iovss.n3358 iovss.n3357 0.00281579
R14461 iovss.n3357 iovss.n3356 0.00281579
R14462 iovss.n3356 iovss.n3355 0.00281579
R14463 iovss.n3355 iovss.n3354 0.00281579
R14464 iovss.n3354 iovss.n3353 0.00281579
R14465 iovss.n3353 iovss.n3352 0.00281579
R14466 iovss.n3352 iovss.n3351 0.00281579
R14467 iovss.n3351 iovss.n3350 0.00281579
R14468 iovss.n3350 iovss.n3349 0.00281579
R14469 iovss.n3349 iovss.n3348 0.00281579
R14470 iovss.n3348 iovss.n3347 0.00281579
R14471 iovss.n3347 iovss.n3346 0.00281579
R14472 iovss.n3346 iovss.n3345 0.00281579
R14473 iovss.n3345 iovss.n264 0.00281579
R14474 iovss.n3395 iovss.n264 0.00281579
R14475 iovss.n3413 iovss.n3412 0.00281579
R14476 iovss.n3412 iovss.n3411 0.00281579
R14477 iovss.n3411 iovss.n3410 0.00281579
R14478 iovss.n3410 iovss.n3409 0.00281579
R14479 iovss.n3409 iovss.n3408 0.00281579
R14480 iovss.n3408 iovss.n3407 0.00281579
R14481 iovss.n3407 iovss.n3406 0.00281579
R14482 iovss.n3406 iovss.n3405 0.00281579
R14483 iovss.n3405 iovss.n3404 0.00281579
R14484 iovss.n3404 iovss.n3403 0.00281579
R14485 iovss.n3403 iovss.n3402 0.00281579
R14486 iovss.n3402 iovss.n3401 0.00281579
R14487 iovss.n3401 iovss.n3400 0.00281579
R14488 iovss.n3400 iovss.n3399 0.00281579
R14489 iovss.n3399 iovss.n3398 0.00281579
R14490 iovss.n3398 iovss.n3397 0.00281579
R14491 iovss.n3397 iovss.n3396 0.00281579
R14492 iovss.n3396 iovss.n173 0.00281579
R14493 iovss.n3430 iovss.n174 0.00281579
R14494 iovss.n1321 iovss.n174 0.00281579
R14495 iovss.n1322 iovss.n1321 0.00281579
R14496 iovss.n1323 iovss.n1322 0.00281579
R14497 iovss.n1324 iovss.n1323 0.00281579
R14498 iovss.n1325 iovss.n1324 0.00281579
R14499 iovss.n1326 iovss.n1325 0.00281579
R14500 iovss.n1327 iovss.n1326 0.00281579
R14501 iovss.n1328 iovss.n1327 0.00281579
R14502 iovss.n1329 iovss.n1328 0.00281579
R14503 iovss.n1330 iovss.n1329 0.00281579
R14504 iovss.n1331 iovss.n1330 0.00281579
R14505 iovss.n1332 iovss.n1331 0.00281579
R14506 iovss.n1333 iovss.n1332 0.00281579
R14507 iovss.n1334 iovss.n1333 0.00281579
R14508 iovss.n1335 iovss.n1334 0.00281579
R14509 iovss.n1336 iovss.n1335 0.00281579
R14510 iovss.n1337 iovss.n1336 0.00281579
R14511 iovss.n3437 iovss.n78 0.0027
R14512 iovss.n1137 iovss.n1114 0.00261959
R14513 iovss.n883 iovss 0.00261765
R14514 iovss.n2067 iovss.n2028 0.00255333
R14515 iovss.n2587 iovss.n1434 0.00255333
R14516 iovss.n3103 iovss.n3102 0.00248367
R14517 iovss.n3339 iovss.n3338 0.00248
R14518 iovss.n3465 iovss.n55 0.002425
R14519 iovss.n2753 iovss.n1116 0.00239804
R14520 iovss.n2760 iovss.n876 0.00239804
R14521 iovss.n3260 iovss.n489 0.00237
R14522 iovss.n144 iovss.n105 0.00226
R14523 iovss.n46 iovss.n45 0.00224473
R14524 iovss.n2241 iovss.n2240 0.00219098
R14525 iovss.n2751 iovss.n2602 0.00219098
R14526 iovss.n2886 iovss.n1219 0.00219098
R14527 iovss.n3390 iovss.n358 0.00219098
R14528 iovss.n3427 iovss.n263 0.00219098
R14529 iovss.n263 iovss.n253 0.00219098
R14530 iovss.n949 iovss.n930 0.00219098
R14531 iovss.n3130 iovss.n930 0.00219098
R14532 iovss.n2760 iovss.n1341 0.00219098
R14533 iovss.n1198 iovss.n907 0.00219098
R14534 iovss.n1312 iovss.n1309 0.00219098
R14535 iovss.n3144 iovss.n886 0.00219098
R14536 iovss.n3435 iovss.n119 0.00216715
R14537 iovss.n164 iovss.n93 0.00216715
R14538 iovss.n165 iovss.n92 0.00216715
R14539 iovss.n166 iovss.n91 0.00216715
R14540 iovss.n167 iovss.n90 0.00216715
R14541 iovss.n168 iovss.n89 0.00216715
R14542 iovss.n169 iovss.n88 0.00216715
R14543 iovss.n169 iovss.n85 0.00216715
R14544 iovss.n168 iovss.n84 0.00216715
R14545 iovss.n167 iovss.n83 0.00216715
R14546 iovss.n166 iovss.n82 0.00216715
R14547 iovss.n165 iovss.n81 0.00216715
R14548 iovss.n164 iovss.n80 0.00216715
R14549 iovss.n119 iovss.n79 0.00216715
R14550 iovss.n2393 iovss.n2356 0.00216715
R14551 iovss.n1676 iovss.n1627 0.00216715
R14552 iovss.n1675 iovss.n1628 0.00216715
R14553 iovss.n1674 iovss.n1629 0.00216715
R14554 iovss.n1673 iovss.n1630 0.00216715
R14555 iovss.n1672 iovss.n1631 0.00216715
R14556 iovss.n1671 iovss.n1632 0.00216715
R14557 iovss.n1670 iovss.n1633 0.00216715
R14558 iovss.n1669 iovss.n1634 0.00216715
R14559 iovss.n1668 iovss.n1635 0.00216715
R14560 iovss.n1667 iovss.n1636 0.00216715
R14561 iovss.n1666 iovss.n1637 0.00216715
R14562 iovss.n1665 iovss.n1638 0.00216715
R14563 iovss.n1664 iovss.n1639 0.00216715
R14564 iovss.n1663 iovss.n1640 0.00216715
R14565 iovss.n1662 iovss.n1641 0.00216715
R14566 iovss.n1661 iovss.n1642 0.00216715
R14567 iovss.n1660 iovss.n1643 0.00216715
R14568 iovss.n1659 iovss.n1644 0.00216715
R14569 iovss.n1658 iovss.n1645 0.00216715
R14570 iovss.n1657 iovss.n1646 0.00216715
R14571 iovss.n1656 iovss.n1647 0.00216715
R14572 iovss.n1655 iovss.n1648 0.00216715
R14573 iovss.n1654 iovss.n1649 0.00216715
R14574 iovss.n2395 iovss.n1650 0.00216715
R14575 iovss.n2397 iovss.n1549 0.00216715
R14576 iovss.n2356 iovss.n220 0.00216715
R14577 iovss.n1676 iovss.n1624 0.00216715
R14578 iovss.n1675 iovss.n1623 0.00216715
R14579 iovss.n1674 iovss.n1622 0.00216715
R14580 iovss.n1673 iovss.n1621 0.00216715
R14581 iovss.n1672 iovss.n1620 0.00216715
R14582 iovss.n1671 iovss.n1619 0.00216715
R14583 iovss.n1670 iovss.n1618 0.00216715
R14584 iovss.n1669 iovss.n1617 0.00216715
R14585 iovss.n1668 iovss.n1616 0.00216715
R14586 iovss.n1667 iovss.n1615 0.00216715
R14587 iovss.n1666 iovss.n1614 0.00216715
R14588 iovss.n1665 iovss.n1613 0.00216715
R14589 iovss.n1664 iovss.n1612 0.00216715
R14590 iovss.n1663 iovss.n1611 0.00216715
R14591 iovss.n1662 iovss.n1610 0.00216715
R14592 iovss.n1661 iovss.n1609 0.00216715
R14593 iovss.n1660 iovss.n1608 0.00216715
R14594 iovss.n1659 iovss.n1607 0.00216715
R14595 iovss.n1658 iovss.n1606 0.00216715
R14596 iovss.n1657 iovss.n1605 0.00216715
R14597 iovss.n1656 iovss.n1604 0.00216715
R14598 iovss.n1655 iovss.n1603 0.00216715
R14599 iovss.n1654 iovss.n1602 0.00216715
R14600 iovss.n1650 iovss.n1601 0.00216715
R14601 iovss.n1600 iovss.n1549 0.00216715
R14602 iovss.n733 iovss.n646 0.00216715
R14603 iovss.n765 iovss.n644 0.00216715
R14604 iovss.n734 iovss.n647 0.00216715
R14605 iovss.n764 iovss.n643 0.00216715
R14606 iovss.n735 iovss.n648 0.00216715
R14607 iovss.n763 iovss.n642 0.00216715
R14608 iovss.n736 iovss.n649 0.00216715
R14609 iovss.n762 iovss.n641 0.00216715
R14610 iovss.n737 iovss.n650 0.00216715
R14611 iovss.n761 iovss.n640 0.00216715
R14612 iovss.n738 iovss.n651 0.00216715
R14613 iovss.n760 iovss.n639 0.00216715
R14614 iovss.n739 iovss.n652 0.00216715
R14615 iovss.n759 iovss.n638 0.00216715
R14616 iovss.n740 iovss.n653 0.00216715
R14617 iovss.n758 iovss.n637 0.00216715
R14618 iovss.n741 iovss.n654 0.00216715
R14619 iovss.n757 iovss.n636 0.00216715
R14620 iovss.n3250 iovss.n655 0.00216715
R14621 iovss.n2215 iovss.n1918 0.00216715
R14622 iovss.n2156 iovss.n1916 0.00216715
R14623 iovss.n2216 iovss.n1919 0.00216715
R14624 iovss.n2155 iovss.n1915 0.00216715
R14625 iovss.n2217 iovss.n1920 0.00216715
R14626 iovss.n2154 iovss.n1914 0.00216715
R14627 iovss.n2218 iovss.n1921 0.00216715
R14628 iovss.n2153 iovss.n1913 0.00216715
R14629 iovss.n2219 iovss.n1922 0.00216715
R14630 iovss.n2152 iovss.n1912 0.00216715
R14631 iovss.n2220 iovss.n1923 0.00216715
R14632 iovss.n2151 iovss.n1911 0.00216715
R14633 iovss.n2221 iovss.n1924 0.00216715
R14634 iovss.n2150 iovss.n1910 0.00216715
R14635 iovss.n2222 iovss.n1925 0.00216715
R14636 iovss.n2149 iovss.n1909 0.00216715
R14637 iovss.n2223 iovss.n1926 0.00216715
R14638 iovss.n2148 iovss.n1908 0.00216715
R14639 iovss.n2224 iovss.n1927 0.00216715
R14640 iovss.n2147 iovss.n1907 0.00216715
R14641 iovss.n2225 iovss.n1928 0.00216715
R14642 iovss.n2146 iovss.n1906 0.00216715
R14643 iovss.n2226 iovss.n1929 0.00216715
R14644 iovss.n2145 iovss.n1905 0.00216715
R14645 iovss.n2227 iovss.n1930 0.00216715
R14646 iovss.n2144 iovss.n1904 0.00216715
R14647 iovss.n2228 iovss.n1931 0.00216715
R14648 iovss.n2143 iovss.n1903 0.00216715
R14649 iovss.n2229 iovss.n1932 0.00216715
R14650 iovss.n2142 iovss.n1902 0.00216715
R14651 iovss.n2230 iovss.n1933 0.00216715
R14652 iovss.n2141 iovss.n1901 0.00216715
R14653 iovss.n2231 iovss.n1934 0.00216715
R14654 iovss.n2140 iovss.n1900 0.00216715
R14655 iovss.n2232 iovss.n1935 0.00216715
R14656 iovss.n2139 iovss.n1899 0.00216715
R14657 iovss.n2233 iovss.n1936 0.00216715
R14658 iovss.n2138 iovss.n1898 0.00216715
R14659 iovss.n2234 iovss.n1937 0.00216715
R14660 iovss.n2137 iovss.n1897 0.00216715
R14661 iovss.n2235 iovss.n1938 0.00216715
R14662 iovss.n2136 iovss.n1896 0.00216715
R14663 iovss.n2236 iovss.n1939 0.00216715
R14664 iovss.n2135 iovss.n1895 0.00216715
R14665 iovss.n2237 iovss.n1940 0.00216715
R14666 iovss.n2134 iovss.n1894 0.00216715
R14667 iovss.n2238 iovss.n1941 0.00216715
R14668 iovss.n2133 iovss.n1893 0.00216715
R14669 iovss.n2239 iovss.n1942 0.00216715
R14670 iovss.n2132 iovss.n1892 0.00216715
R14671 iovss.n2242 iovss.n1943 0.00216715
R14672 iovss.n2089 iovss.n1973 0.00216715
R14673 iovss.n2079 iovss.n1440 0.00216715
R14674 iovss.n1998 iovss.n1982 0.00216715
R14675 iovss.n2091 iovss.n1997 0.00216715
R14676 iovss.n2093 iovss.n1973 0.00216715
R14677 iovss.n2089 iovss.n2079 0.00216715
R14678 iovss.n1998 iovss.n1441 0.00216715
R14679 iovss.n1997 iovss.n1982 0.00216715
R14680 iovss.n3391 iovss.n335 0.00216715
R14681 iovss.n336 iovss.n274 0.00216715
R14682 iovss.n350 iovss.n277 0.00216715
R14683 iovss.n3385 iovss.n273 0.00216715
R14684 iovss.n351 iovss.n278 0.00216715
R14685 iovss.n3384 iovss.n272 0.00216715
R14686 iovss.n352 iovss.n279 0.00216715
R14687 iovss.n3383 iovss.n271 0.00216715
R14688 iovss.n353 iovss.n280 0.00216715
R14689 iovss.n3382 iovss.n270 0.00216715
R14690 iovss.n354 iovss.n281 0.00216715
R14691 iovss.n3381 iovss.n269 0.00216715
R14692 iovss.n355 iovss.n282 0.00216715
R14693 iovss.n3380 iovss.n268 0.00216715
R14694 iovss.n356 iovss.n283 0.00216715
R14695 iovss.n3379 iovss.n267 0.00216715
R14696 iovss.n357 iovss.n284 0.00216715
R14697 iovss.n3378 iovss.n266 0.00216715
R14698 iovss.n3393 iovss.n285 0.00216715
R14699 iovss.n2289 iovss.n1732 0.00216715
R14700 iovss.n1782 iovss.n1730 0.00216715
R14701 iovss.n1844 iovss.n1733 0.00216715
R14702 iovss.n1781 iovss.n1729 0.00216715
R14703 iovss.n1845 iovss.n1734 0.00216715
R14704 iovss.n1780 iovss.n1728 0.00216715
R14705 iovss.n1846 iovss.n1735 0.00216715
R14706 iovss.n1779 iovss.n1727 0.00216715
R14707 iovss.n1847 iovss.n1736 0.00216715
R14708 iovss.n1778 iovss.n1726 0.00216715
R14709 iovss.n1848 iovss.n1737 0.00216715
R14710 iovss.n1777 iovss.n1725 0.00216715
R14711 iovss.n1849 iovss.n1738 0.00216715
R14712 iovss.n1776 iovss.n1724 0.00216715
R14713 iovss.n1850 iovss.n1739 0.00216715
R14714 iovss.n1775 iovss.n1723 0.00216715
R14715 iovss.n1851 iovss.n1740 0.00216715
R14716 iovss.n1774 iovss.n1722 0.00216715
R14717 iovss.n1852 iovss.n1741 0.00216715
R14718 iovss.n1773 iovss.n1721 0.00216715
R14719 iovss.n1853 iovss.n1742 0.00216715
R14720 iovss.n1772 iovss.n1720 0.00216715
R14721 iovss.n1854 iovss.n1743 0.00216715
R14722 iovss.n1771 iovss.n1719 0.00216715
R14723 iovss.n1855 iovss.n1744 0.00216715
R14724 iovss.n1770 iovss.n1718 0.00216715
R14725 iovss.n1856 iovss.n1745 0.00216715
R14726 iovss.n1769 iovss.n1717 0.00216715
R14727 iovss.n1857 iovss.n1746 0.00216715
R14728 iovss.n1768 iovss.n1716 0.00216715
R14729 iovss.n1858 iovss.n1747 0.00216715
R14730 iovss.n1767 iovss.n1715 0.00216715
R14731 iovss.n1859 iovss.n1748 0.00216715
R14732 iovss.n1766 iovss.n1714 0.00216715
R14733 iovss.n1860 iovss.n1749 0.00216715
R14734 iovss.n1765 iovss.n1713 0.00216715
R14735 iovss.n1861 iovss.n1750 0.00216715
R14736 iovss.n1764 iovss.n1712 0.00216715
R14737 iovss.n1862 iovss.n1751 0.00216715
R14738 iovss.n1763 iovss.n1711 0.00216715
R14739 iovss.n1863 iovss.n1752 0.00216715
R14740 iovss.n1762 iovss.n1710 0.00216715
R14741 iovss.n1864 iovss.n1753 0.00216715
R14742 iovss.n1761 iovss.n1709 0.00216715
R14743 iovss.n1865 iovss.n1754 0.00216715
R14744 iovss.n1760 iovss.n1708 0.00216715
R14745 iovss.n1866 iovss.n1755 0.00216715
R14746 iovss.n1759 iovss.n1707 0.00216715
R14747 iovss.n1867 iovss.n1756 0.00216715
R14748 iovss.n1758 iovss.n1706 0.00216715
R14749 iovss.n2291 iovss.n1757 0.00216715
R14750 iovss.n2557 iovss.n2552 0.00216715
R14751 iovss.n2553 iovss.n1448 0.00216715
R14752 iovss.n1486 iovss.n1449 0.00216715
R14753 iovss.n2561 iovss.n2556 0.00216715
R14754 iovss.n2557 iovss.n1502 0.00216715
R14755 iovss.n2553 iovss.n2552 0.00216715
R14756 iovss.n2563 iovss.n1449 0.00216715
R14757 iovss.n2556 iovss.n1486 0.00216715
R14758 iovss.n2289 iovss.n303 0.00216715
R14759 iovss.n1782 iovss.n1732 0.00216715
R14760 iovss.n1844 iovss.n1730 0.00216715
R14761 iovss.n1781 iovss.n1733 0.00216715
R14762 iovss.n1845 iovss.n1729 0.00216715
R14763 iovss.n1780 iovss.n1734 0.00216715
R14764 iovss.n1846 iovss.n1728 0.00216715
R14765 iovss.n1779 iovss.n1735 0.00216715
R14766 iovss.n1847 iovss.n1727 0.00216715
R14767 iovss.n1778 iovss.n1736 0.00216715
R14768 iovss.n1848 iovss.n1726 0.00216715
R14769 iovss.n1777 iovss.n1737 0.00216715
R14770 iovss.n1849 iovss.n1725 0.00216715
R14771 iovss.n1776 iovss.n1738 0.00216715
R14772 iovss.n1850 iovss.n1724 0.00216715
R14773 iovss.n1775 iovss.n1739 0.00216715
R14774 iovss.n1851 iovss.n1723 0.00216715
R14775 iovss.n1774 iovss.n1740 0.00216715
R14776 iovss.n1852 iovss.n1722 0.00216715
R14777 iovss.n1773 iovss.n1741 0.00216715
R14778 iovss.n1853 iovss.n1721 0.00216715
R14779 iovss.n1772 iovss.n1742 0.00216715
R14780 iovss.n1854 iovss.n1720 0.00216715
R14781 iovss.n1771 iovss.n1743 0.00216715
R14782 iovss.n1855 iovss.n1719 0.00216715
R14783 iovss.n1770 iovss.n1744 0.00216715
R14784 iovss.n1856 iovss.n1718 0.00216715
R14785 iovss.n1769 iovss.n1745 0.00216715
R14786 iovss.n1857 iovss.n1717 0.00216715
R14787 iovss.n1768 iovss.n1746 0.00216715
R14788 iovss.n1858 iovss.n1716 0.00216715
R14789 iovss.n1767 iovss.n1747 0.00216715
R14790 iovss.n1859 iovss.n1715 0.00216715
R14791 iovss.n1766 iovss.n1748 0.00216715
R14792 iovss.n1860 iovss.n1714 0.00216715
R14793 iovss.n1765 iovss.n1749 0.00216715
R14794 iovss.n1861 iovss.n1713 0.00216715
R14795 iovss.n1764 iovss.n1750 0.00216715
R14796 iovss.n1862 iovss.n1712 0.00216715
R14797 iovss.n1763 iovss.n1751 0.00216715
R14798 iovss.n1863 iovss.n1711 0.00216715
R14799 iovss.n1762 iovss.n1752 0.00216715
R14800 iovss.n1864 iovss.n1710 0.00216715
R14801 iovss.n1761 iovss.n1753 0.00216715
R14802 iovss.n1865 iovss.n1709 0.00216715
R14803 iovss.n1760 iovss.n1754 0.00216715
R14804 iovss.n1866 iovss.n1708 0.00216715
R14805 iovss.n1759 iovss.n1755 0.00216715
R14806 iovss.n1867 iovss.n1707 0.00216715
R14807 iovss.n1758 iovss.n1756 0.00216715
R14808 iovss.n1757 iovss.n1706 0.00216715
R14809 iovss.n2215 iovss.n673 0.00216715
R14810 iovss.n2156 iovss.n1918 0.00216715
R14811 iovss.n2216 iovss.n1916 0.00216715
R14812 iovss.n2155 iovss.n1919 0.00216715
R14813 iovss.n2217 iovss.n1915 0.00216715
R14814 iovss.n2154 iovss.n1920 0.00216715
R14815 iovss.n2218 iovss.n1914 0.00216715
R14816 iovss.n2153 iovss.n1921 0.00216715
R14817 iovss.n2219 iovss.n1913 0.00216715
R14818 iovss.n2152 iovss.n1922 0.00216715
R14819 iovss.n2220 iovss.n1912 0.00216715
R14820 iovss.n2151 iovss.n1923 0.00216715
R14821 iovss.n2221 iovss.n1911 0.00216715
R14822 iovss.n2150 iovss.n1924 0.00216715
R14823 iovss.n2222 iovss.n1910 0.00216715
R14824 iovss.n2149 iovss.n1925 0.00216715
R14825 iovss.n2223 iovss.n1909 0.00216715
R14826 iovss.n2148 iovss.n1926 0.00216715
R14827 iovss.n2224 iovss.n1908 0.00216715
R14828 iovss.n2147 iovss.n1927 0.00216715
R14829 iovss.n2225 iovss.n1907 0.00216715
R14830 iovss.n2146 iovss.n1928 0.00216715
R14831 iovss.n2226 iovss.n1906 0.00216715
R14832 iovss.n2145 iovss.n1929 0.00216715
R14833 iovss.n2227 iovss.n1905 0.00216715
R14834 iovss.n2144 iovss.n1930 0.00216715
R14835 iovss.n2228 iovss.n1904 0.00216715
R14836 iovss.n2143 iovss.n1931 0.00216715
R14837 iovss.n2229 iovss.n1903 0.00216715
R14838 iovss.n2142 iovss.n1932 0.00216715
R14839 iovss.n2230 iovss.n1902 0.00216715
R14840 iovss.n2141 iovss.n1933 0.00216715
R14841 iovss.n2231 iovss.n1901 0.00216715
R14842 iovss.n2140 iovss.n1934 0.00216715
R14843 iovss.n2232 iovss.n1900 0.00216715
R14844 iovss.n2139 iovss.n1935 0.00216715
R14845 iovss.n2233 iovss.n1899 0.00216715
R14846 iovss.n2138 iovss.n1936 0.00216715
R14847 iovss.n2234 iovss.n1898 0.00216715
R14848 iovss.n2137 iovss.n1937 0.00216715
R14849 iovss.n2235 iovss.n1897 0.00216715
R14850 iovss.n2136 iovss.n1938 0.00216715
R14851 iovss.n2236 iovss.n1896 0.00216715
R14852 iovss.n2135 iovss.n1939 0.00216715
R14853 iovss.n2237 iovss.n1895 0.00216715
R14854 iovss.n2134 iovss.n1940 0.00216715
R14855 iovss.n2238 iovss.n1894 0.00216715
R14856 iovss.n2133 iovss.n1941 0.00216715
R14857 iovss.n2239 iovss.n1893 0.00216715
R14858 iovss.n2132 iovss.n1942 0.00216715
R14859 iovss.n1943 iovss.n1892 0.00216715
R14860 iovss.n411 iovss.n381 0.00216715
R14861 iovss.n408 iovss.n401 0.00216715
R14862 iovss.n400 iovss.n382 0.00216715
R14863 iovss.n407 iovss.n399 0.00216715
R14864 iovss.n398 iovss.n383 0.00216715
R14865 iovss.n406 iovss.n397 0.00216715
R14866 iovss.n396 iovss.n384 0.00216715
R14867 iovss.n405 iovss.n395 0.00216715
R14868 iovss.n394 iovss.n385 0.00216715
R14869 iovss.n404 iovss.n393 0.00216715
R14870 iovss.n392 iovss.n386 0.00216715
R14871 iovss.n403 iovss.n391 0.00216715
R14872 iovss.n390 iovss.n387 0.00216715
R14873 iovss.n402 iovss.n389 0.00216715
R14874 iovss.n3344 iovss.n360 0.00216715
R14875 iovss.n520 iovss.n490 0.00216715
R14876 iovss.n517 iovss.n510 0.00216715
R14877 iovss.n509 iovss.n491 0.00216715
R14878 iovss.n516 iovss.n508 0.00216715
R14879 iovss.n507 iovss.n492 0.00216715
R14880 iovss.n515 iovss.n506 0.00216715
R14881 iovss.n505 iovss.n493 0.00216715
R14882 iovss.n514 iovss.n504 0.00216715
R14883 iovss.n503 iovss.n494 0.00216715
R14884 iovss.n513 iovss.n502 0.00216715
R14885 iovss.n501 iovss.n495 0.00216715
R14886 iovss.n512 iovss.n500 0.00216715
R14887 iovss.n499 iovss.n496 0.00216715
R14888 iovss.n511 iovss.n498 0.00216715
R14889 iovss.n3254 iovss.n615 0.00216715
R14890 iovss.n615 iovss.n498 0.00216715
R14891 iovss.n511 iovss.n496 0.00216715
R14892 iovss.n500 iovss.n499 0.00216715
R14893 iovss.n512 iovss.n495 0.00216715
R14894 iovss.n502 iovss.n501 0.00216715
R14895 iovss.n513 iovss.n494 0.00216715
R14896 iovss.n504 iovss.n503 0.00216715
R14897 iovss.n514 iovss.n493 0.00216715
R14898 iovss.n506 iovss.n505 0.00216715
R14899 iovss.n515 iovss.n492 0.00216715
R14900 iovss.n508 iovss.n507 0.00216715
R14901 iovss.n516 iovss.n491 0.00216715
R14902 iovss.n510 iovss.n509 0.00216715
R14903 iovss.n517 iovss.n490 0.00216715
R14904 iovss.n3258 iovss.n520 0.00216715
R14905 iovss.n389 iovss.n360 0.00216715
R14906 iovss.n402 iovss.n387 0.00216715
R14907 iovss.n391 iovss.n390 0.00216715
R14908 iovss.n403 iovss.n386 0.00216715
R14909 iovss.n393 iovss.n392 0.00216715
R14910 iovss.n404 iovss.n385 0.00216715
R14911 iovss.n395 iovss.n394 0.00216715
R14912 iovss.n405 iovss.n384 0.00216715
R14913 iovss.n397 iovss.n396 0.00216715
R14914 iovss.n406 iovss.n383 0.00216715
R14915 iovss.n399 iovss.n398 0.00216715
R14916 iovss.n407 iovss.n382 0.00216715
R14917 iovss.n401 iovss.n400 0.00216715
R14918 iovss.n408 iovss.n381 0.00216715
R14919 iovss.n3342 iovss.n411 0.00216715
R14920 iovss.n100 iovss.n93 0.00216715
R14921 iovss.n99 iovss.n92 0.00216715
R14922 iovss.n98 iovss.n91 0.00216715
R14923 iovss.n97 iovss.n90 0.00216715
R14924 iovss.n96 iovss.n89 0.00216715
R14925 iovss.n95 iovss.n88 0.00216715
R14926 iovss.n102 iovss.n87 0.00216715
R14927 iovss.n3432 iovss.n149 0.00216715
R14928 iovss.n149 iovss.n87 0.00216715
R14929 iovss.n102 iovss.n85 0.00216715
R14930 iovss.n95 iovss.n84 0.00216715
R14931 iovss.n96 iovss.n83 0.00216715
R14932 iovss.n97 iovss.n82 0.00216715
R14933 iovss.n98 iovss.n81 0.00216715
R14934 iovss.n99 iovss.n80 0.00216715
R14935 iovss.n100 iovss.n79 0.00216715
R14936 iovss.n3426 iovss.n3414 0.00216715
R14937 iovss.n3415 iovss.n184 0.00216715
R14938 iovss.n255 iovss.n186 0.00216715
R14939 iovss.n202 iovss.n183 0.00216715
R14940 iovss.n256 iovss.n187 0.00216715
R14941 iovss.n201 iovss.n182 0.00216715
R14942 iovss.n257 iovss.n188 0.00216715
R14943 iovss.n200 iovss.n181 0.00216715
R14944 iovss.n258 iovss.n189 0.00216715
R14945 iovss.n199 iovss.n180 0.00216715
R14946 iovss.n259 iovss.n190 0.00216715
R14947 iovss.n198 iovss.n179 0.00216715
R14948 iovss.n260 iovss.n191 0.00216715
R14949 iovss.n197 iovss.n178 0.00216715
R14950 iovss.n261 iovss.n192 0.00216715
R14951 iovss.n196 iovss.n177 0.00216715
R14952 iovss.n262 iovss.n193 0.00216715
R14953 iovss.n195 iovss.n176 0.00216715
R14954 iovss.n3428 iovss.n194 0.00216715
R14955 iovss.n2381 iovss.n1624 0.00216715
R14956 iovss.n2379 iovss.n1623 0.00216715
R14957 iovss.n2378 iovss.n1622 0.00216715
R14958 iovss.n2377 iovss.n1621 0.00216715
R14959 iovss.n2376 iovss.n1620 0.00216715
R14960 iovss.n2375 iovss.n1619 0.00216715
R14961 iovss.n2374 iovss.n1618 0.00216715
R14962 iovss.n2373 iovss.n1617 0.00216715
R14963 iovss.n2372 iovss.n1616 0.00216715
R14964 iovss.n2371 iovss.n1615 0.00216715
R14965 iovss.n2370 iovss.n1614 0.00216715
R14966 iovss.n2369 iovss.n1613 0.00216715
R14967 iovss.n2368 iovss.n1612 0.00216715
R14968 iovss.n2367 iovss.n1611 0.00216715
R14969 iovss.n2366 iovss.n1610 0.00216715
R14970 iovss.n2365 iovss.n1609 0.00216715
R14971 iovss.n2364 iovss.n1608 0.00216715
R14972 iovss.n2363 iovss.n1607 0.00216715
R14973 iovss.n2362 iovss.n1606 0.00216715
R14974 iovss.n2361 iovss.n1605 0.00216715
R14975 iovss.n2360 iovss.n1604 0.00216715
R14976 iovss.n2359 iovss.n1603 0.00216715
R14977 iovss.n2358 iovss.n1602 0.00216715
R14978 iovss.n2357 iovss.n1601 0.00216715
R14979 iovss.n1651 iovss.n1600 0.00216715
R14980 iovss.n2507 iovss.n2399 0.00216715
R14981 iovss.n2402 iovss.n1444 0.00216715
R14982 iovss.n2401 iovss.n1548 0.00216715
R14983 iovss.n2502 iovss.n2400 0.00216715
R14984 iovss.n2393 iovss.n2381 0.00216715
R14985 iovss.n2379 iovss.n1627 0.00216715
R14986 iovss.n2378 iovss.n1628 0.00216715
R14987 iovss.n2377 iovss.n1629 0.00216715
R14988 iovss.n2376 iovss.n1630 0.00216715
R14989 iovss.n2375 iovss.n1631 0.00216715
R14990 iovss.n2374 iovss.n1632 0.00216715
R14991 iovss.n2373 iovss.n1633 0.00216715
R14992 iovss.n2372 iovss.n1634 0.00216715
R14993 iovss.n2371 iovss.n1635 0.00216715
R14994 iovss.n2370 iovss.n1636 0.00216715
R14995 iovss.n2369 iovss.n1637 0.00216715
R14996 iovss.n2368 iovss.n1638 0.00216715
R14997 iovss.n2367 iovss.n1639 0.00216715
R14998 iovss.n2366 iovss.n1640 0.00216715
R14999 iovss.n2365 iovss.n1641 0.00216715
R15000 iovss.n2364 iovss.n1642 0.00216715
R15001 iovss.n2363 iovss.n1643 0.00216715
R15002 iovss.n2362 iovss.n1644 0.00216715
R15003 iovss.n2361 iovss.n1645 0.00216715
R15004 iovss.n2360 iovss.n1646 0.00216715
R15005 iovss.n2359 iovss.n1647 0.00216715
R15006 iovss.n2358 iovss.n1648 0.00216715
R15007 iovss.n2357 iovss.n1649 0.00216715
R15008 iovss.n2395 iovss.n1651 0.00216715
R15009 iovss.n2507 iovss.n2398 0.00216715
R15010 iovss.n2402 iovss.n2399 0.00216715
R15011 iovss.n2401 iovss.n1443 0.00216715
R15012 iovss.n2502 iovss.n1548 0.00216715
R15013 iovss.n3414 iovss.n172 0.00216715
R15014 iovss.n3426 iovss.n3415 0.00216715
R15015 iovss.n255 iovss.n184 0.00216715
R15016 iovss.n202 iovss.n186 0.00216715
R15017 iovss.n256 iovss.n183 0.00216715
R15018 iovss.n201 iovss.n187 0.00216715
R15019 iovss.n257 iovss.n182 0.00216715
R15020 iovss.n200 iovss.n188 0.00216715
R15021 iovss.n258 iovss.n181 0.00216715
R15022 iovss.n199 iovss.n189 0.00216715
R15023 iovss.n259 iovss.n180 0.00216715
R15024 iovss.n198 iovss.n190 0.00216715
R15025 iovss.n260 iovss.n179 0.00216715
R15026 iovss.n197 iovss.n191 0.00216715
R15027 iovss.n261 iovss.n178 0.00216715
R15028 iovss.n196 iovss.n192 0.00216715
R15029 iovss.n262 iovss.n177 0.00216715
R15030 iovss.n195 iovss.n193 0.00216715
R15031 iovss.n194 iovss.n176 0.00216715
R15032 iovss.n335 iovss.n275 0.00216715
R15033 iovss.n3391 iovss.n336 0.00216715
R15034 iovss.n350 iovss.n274 0.00216715
R15035 iovss.n3385 iovss.n277 0.00216715
R15036 iovss.n351 iovss.n273 0.00216715
R15037 iovss.n3384 iovss.n278 0.00216715
R15038 iovss.n352 iovss.n272 0.00216715
R15039 iovss.n3383 iovss.n279 0.00216715
R15040 iovss.n353 iovss.n271 0.00216715
R15041 iovss.n3382 iovss.n280 0.00216715
R15042 iovss.n354 iovss.n270 0.00216715
R15043 iovss.n3381 iovss.n281 0.00216715
R15044 iovss.n355 iovss.n269 0.00216715
R15045 iovss.n3380 iovss.n282 0.00216715
R15046 iovss.n356 iovss.n268 0.00216715
R15047 iovss.n3379 iovss.n283 0.00216715
R15048 iovss.n357 iovss.n267 0.00216715
R15049 iovss.n3378 iovss.n284 0.00216715
R15050 iovss.n285 iovss.n266 0.00216715
R15051 iovss.n733 iovss.n632 0.00216715
R15052 iovss.n765 iovss.n646 0.00216715
R15053 iovss.n734 iovss.n644 0.00216715
R15054 iovss.n764 iovss.n647 0.00216715
R15055 iovss.n735 iovss.n643 0.00216715
R15056 iovss.n763 iovss.n648 0.00216715
R15057 iovss.n736 iovss.n642 0.00216715
R15058 iovss.n762 iovss.n649 0.00216715
R15059 iovss.n737 iovss.n641 0.00216715
R15060 iovss.n761 iovss.n650 0.00216715
R15061 iovss.n738 iovss.n640 0.00216715
R15062 iovss.n760 iovss.n651 0.00216715
R15063 iovss.n739 iovss.n639 0.00216715
R15064 iovss.n759 iovss.n652 0.00216715
R15065 iovss.n740 iovss.n638 0.00216715
R15066 iovss.n758 iovss.n653 0.00216715
R15067 iovss.n741 iovss.n637 0.00216715
R15068 iovss.n757 iovss.n654 0.00216715
R15069 iovss.n655 iovss.n636 0.00216715
R15070 iovss.n2205 iovss.n1952 0.00215647
R15071 iovss.n3251 iovss.n635 0.00215647
R15072 iovss.n580 iovss.n536 0.00215
R15073 iovss.n2281 iovss.n1832 0.00212196
R15074 iovss.n2279 iovss.n1824 0.00212196
R15075 iovss.n2602 iovss.n989 0.00212196
R15076 iovss.n811 iovss.n324 0.00212196
R15077 iovss.n819 iovss.n318 0.00212196
R15078 iovss.n1340 iovss.n875 0.00212196
R15079 iovss.n2207 iovss.n1949 0.00208745
R15080 iovss.n783 iovss.n661 0.00208745
R15081 iovss.n1695 iovss.n1553 0.00205294
R15082 iovss.n2309 iovss.n1558 0.00205294
R15083 iovss.n839 iovss.n205 0.00205294
R15084 iovss.n847 iovss.n210 0.00205294
R15085 iovss.n429 iovss.n388 0.00204
R15086 iovss.n452 iovss.n449 0.00204
R15087 iovss.n2203 iovss.n1954 0.00201843
R15088 iovss.n791 iovss.n665 0.00201843
R15089 iovss.n3253 iovss.n632 0.00200081
R15090 iovss.n3362 iovss.n275 0.00200081
R15091 iovss.n3431 iovss.n172 0.00200081
R15092 iovss.n3106 iovss.n3105 0.00199991
R15093 iovss.n2283 iovss.n1837 0.00198392
R15094 iovss.n2277 iovss.n1819 0.00198392
R15095 iovss.n810 iovss.n328 0.00198392
R15096 iovss.n820 iovss.n315 0.00198392
R15097 iovss.n882 iovss 0.00196667
R15098 iovss.n2341 iovss 0.00196667
R15099 iovss.n2043 iovss.n2021 0.00196667
R15100 iovss.n2461 iovss.n2460 0.00196667
R15101 iovss.n2209 iovss.n1947 0.00194941
R15102 iovss.n782 iovss.n659 0.00194941
R15103 iovss.n612 iovss.n522 0.00193
R15104 iovss.n2296 iovss.n1551 0.0019149
R15105 iovss.n2311 iovss.n1560 0.0019149
R15106 iovss.n838 iovss.n203 0.0019149
R15107 iovss.n848 iovss.n211 0.0019149
R15108 iovss.n2182 iovss.n2180 0.00191176
R15109 iovss.n2182 iovss.n2175 0.00191176
R15110 iovss.n2187 iovss.n2175 0.00191176
R15111 iovss.n2189 iovss.n2187 0.00191176
R15112 iovss.n2191 iovss.n2189 0.00191176
R15113 iovss.n2191 iovss.n2172 0.00191176
R15114 iovss.n2198 iovss.n2172 0.00191176
R15115 iovss.n2198 iovss.n2197 0.00191176
R15116 iovss.n2197 iovss.n1887 0.00191176
R15117 iovss.n2250 iovss.n1887 0.00191176
R15118 iovss.n2252 iovss.n2250 0.00191176
R15119 iovss.n2254 iovss.n2252 0.00191176
R15120 iovss.n2254 iovss.n1885 0.00191176
R15121 iovss.n2259 iovss.n1885 0.00191176
R15122 iovss.n2261 iovss.n2259 0.00191176
R15123 iovss.n2263 iovss.n2261 0.00191176
R15124 iovss.n2263 iovss.n1882 0.00191176
R15125 iovss.n2270 iovss.n1882 0.00191176
R15126 iovss.n2270 iovss.n2269 0.00191176
R15127 iovss.n2269 iovss.n1700 0.00191176
R15128 iovss.n2300 iovss.n1700 0.00191176
R15129 iovss.n2300 iovss.n1698 0.00191176
R15130 iovss.n2304 iovss.n1698 0.00191176
R15131 iovss.n2304 iovss.n1692 0.00191176
R15132 iovss.n2315 iovss.n1692 0.00191176
R15133 iovss.n2315 iovss.n1690 0.00191176
R15134 iovss.n2322 iovss.n1690 0.00191176
R15135 iovss.n2322 iovss.n2321 0.00191176
R15136 iovss.n2321 iovss.n1685 0.00191176
R15137 iovss.n2333 iovss.n1685 0.00191176
R15138 iovss.n2335 iovss.n2333 0.00191176
R15139 iovss.n2335 iovss.n1683 0.00191176
R15140 iovss.n2348 iovss.n1683 0.00191176
R15141 iovss.n2348 iovss.n2347 0.00191176
R15142 iovss.n2347 iovss.n2345 0.00191176
R15143 iovss.n2345 iovss.n2343 0.00191176
R15144 iovss.n3241 iovss.n774 0.00191176
R15145 iovss.n3241 iovss.n3240 0.00191176
R15146 iovss.n3240 iovss.n780 0.00191176
R15147 iovss.n3233 iovss.n780 0.00191176
R15148 iovss.n3233 iovss.n3232 0.00191176
R15149 iovss.n3232 iovss.n789 0.00191176
R15150 iovss.n3225 iovss.n789 0.00191176
R15151 iovss.n3225 iovss.n3224 0.00191176
R15152 iovss.n3224 iovss.n799 0.00191176
R15153 iovss.n3217 iovss.n799 0.00191176
R15154 iovss.n3217 iovss.n3216 0.00191176
R15155 iovss.n3216 iovss.n807 0.00191176
R15156 iovss.n3209 iovss.n807 0.00191176
R15157 iovss.n3209 iovss.n3208 0.00191176
R15158 iovss.n3208 iovss.n817 0.00191176
R15159 iovss.n3201 iovss.n817 0.00191176
R15160 iovss.n3201 iovss.n3200 0.00191176
R15161 iovss.n3200 iovss.n827 0.00191176
R15162 iovss.n3193 iovss.n827 0.00191176
R15163 iovss.n3193 iovss.n3192 0.00191176
R15164 iovss.n3192 iovss.n836 0.00191176
R15165 iovss.n3185 iovss.n836 0.00191176
R15166 iovss.n3185 iovss.n3184 0.00191176
R15167 iovss.n3184 iovss.n845 0.00191176
R15168 iovss.n3177 iovss.n845 0.00191176
R15169 iovss.n3177 iovss.n3176 0.00191176
R15170 iovss.n3176 iovss.n854 0.00191176
R15171 iovss.n3169 iovss.n854 0.00191176
R15172 iovss.n3169 iovss.n3168 0.00191176
R15173 iovss.n3168 iovss.n864 0.00191176
R15174 iovss.n3161 iovss.n864 0.00191176
R15175 iovss.n3161 iovss.n3160 0.00191176
R15176 iovss.n3160 iovss.n873 0.00191176
R15177 iovss.n3153 iovss.n873 0.00191176
R15178 iovss.n3153 iovss.n3152 0.00191176
R15179 iovss.n3152 iovss.n883 0.00191176
R15180 iovss.n2721 iovss.n1341 0.00189683
R15181 iovss.n2751 iovss.n2729 0.00189683
R15182 iovss.n2779 iovss.n1309 0.00189683
R15183 iovss.n2886 iovss.n2787 0.00189683
R15184 iovss.n2962 iovss.n886 0.00189683
R15185 iovss.n3070 iovss.n2934 0.00189683
R15186 iovss.n1199 iovss.n1198 0.00189683
R15187 iovss.n1206 iovss.n1115 0.00189683
R15188 iovss.n954 iovss.n930 0.00189683
R15189 iovss.n1056 iovss.n960 0.00189683
R15190 iovss.n2201 iovss.n1956 0.00188039
R15191 iovss.n792 iovss.n667 0.00188039
R15192 iovss.n47 iovss.n46 0.00187364
R15193 iovss.n3249 iovss.n3248 0.00184642
R15194 iovss.n2285 iovss.n1841 0.00184588
R15195 iovss.n2275 iovss.n1814 0.00184588
R15196 iovss.n809 iovss.n331 0.00184588
R15197 iovss.n821 iovss.n312 0.00184588
R15198 iovss.n2157 iovss.n1944 0.00184541
R15199 iovss.n2158 iovss.n2157 0.00184541
R15200 iovss.n2159 iovss.n1945 0.00184541
R15201 iovss.n2130 iovss.n1946 0.00184541
R15202 iovss.n2127 iovss.n1946 0.00184541
R15203 iovss.n2128 iovss.n1947 0.00184541
R15204 iovss.n2125 iovss.n1948 0.00184541
R15205 iovss.n2122 iovss.n1948 0.00184541
R15206 iovss.n2123 iovss.n1949 0.00184541
R15207 iovss.n2120 iovss.n1950 0.00184541
R15208 iovss.n2117 iovss.n1950 0.00184541
R15209 iovss.n2118 iovss.n1951 0.00184541
R15210 iovss.n2115 iovss.n1951 0.00184541
R15211 iovss.n2112 iovss.n1952 0.00184541
R15212 iovss.n2113 iovss.n1953 0.00184541
R15213 iovss.n2110 iovss.n1953 0.00184541
R15214 iovss.n2107 iovss.n1954 0.00184541
R15215 iovss.n2108 iovss.n1955 0.00184541
R15216 iovss.n2105 iovss.n1955 0.00184541
R15217 iovss.n2102 iovss.n1956 0.00184541
R15218 iovss.n2103 iovss.n1957 0.00184541
R15219 iovss.n2099 iovss.n1957 0.00184541
R15220 iovss.n2096 iovss.n1958 0.00184541
R15221 iovss.n2097 iovss.n1960 0.00184541
R15222 iovss.n1960 iovss.n1959 0.00184541
R15223 iovss.n2243 iovss.n1917 0.00184541
R15224 iovss.n2094 iovss.n1961 0.00184541
R15225 iovss.n1842 iovss.n1783 0.00184541
R15226 iovss.n1869 iovss.n1868 0.00184541
R15227 iovss.n1868 iovss.n1843 0.00184541
R15228 iovss.n1838 iovss.n1784 0.00184541
R15229 iovss.n1839 iovss.n1785 0.00184541
R15230 iovss.n1836 iovss.n1785 0.00184541
R15231 iovss.n1833 iovss.n1786 0.00184541
R15232 iovss.n1834 iovss.n1787 0.00184541
R15233 iovss.n1831 iovss.n1787 0.00184541
R15234 iovss.n1828 iovss.n1788 0.00184541
R15235 iovss.n1829 iovss.n1789 0.00184541
R15236 iovss.n1825 iovss.n1789 0.00184541
R15237 iovss.n1826 iovss.n1790 0.00184541
R15238 iovss.n1824 iovss.n1823 0.00184541
R15239 iovss.n1821 iovss.n1791 0.00184541
R15240 iovss.n1822 iovss.n1820 0.00184541
R15241 iovss.n1819 iovss.n1818 0.00184541
R15242 iovss.n1816 iovss.n1793 0.00184541
R15243 iovss.n1817 iovss.n1815 0.00184541
R15244 iovss.n1814 iovss.n1813 0.00184541
R15245 iovss.n1811 iovss.n1795 0.00184541
R15246 iovss.n1812 iovss.n1810 0.00184541
R15247 iovss.n1809 iovss.n1808 0.00184541
R15248 iovss.n1806 iovss.n1797 0.00184541
R15249 iovss.n1807 iovss.n1805 0.00184541
R15250 iovss.n1804 iovss.n1803 0.00184541
R15251 iovss.n1800 iovss.n1799 0.00184541
R15252 iovss.n1801 iovss.n1731 0.00184541
R15253 iovss.n2380 iovss.n1550 0.00184541
R15254 iovss.n2380 iovss.n1625 0.00184541
R15255 iovss.n1626 iovss.n1551 0.00184541
R15256 iovss.n2382 iovss.n1552 0.00184541
R15257 iovss.n1597 iovss.n1552 0.00184541
R15258 iovss.n2383 iovss.n1553 0.00184541
R15259 iovss.n2384 iovss.n1554 0.00184541
R15260 iovss.n1594 iovss.n1554 0.00184541
R15261 iovss.n2385 iovss.n1555 0.00184541
R15262 iovss.n1592 iovss.n1555 0.00184541
R15263 iovss.n2386 iovss.n1556 0.00184541
R15264 iovss.n1590 iovss.n1556 0.00184541
R15265 iovss.n2387 iovss.n1557 0.00184541
R15266 iovss.n1588 iovss.n1557 0.00184541
R15267 iovss.n1586 iovss.n1558 0.00184541
R15268 iovss.n2388 iovss.n1559 0.00184541
R15269 iovss.n1584 iovss.n1559 0.00184541
R15270 iovss.n1582 iovss.n1560 0.00184541
R15271 iovss.n2389 iovss.n1561 0.00184541
R15272 iovss.n1580 iovss.n1561 0.00184541
R15273 iovss.n1578 iovss.n1562 0.00184541
R15274 iovss.n2390 iovss.n1563 0.00184541
R15275 iovss.n1576 iovss.n1563 0.00184541
R15276 iovss.n1574 iovss.n1564 0.00184541
R15277 iovss.n2391 iovss.n1565 0.00184541
R15278 iovss.n1572 iovss.n1565 0.00184541
R15279 iovss.n1570 iovss.n1566 0.00184541
R15280 iovss.n2392 iovss.n1567 0.00184541
R15281 iovss.n1568 iovss.n1567 0.00184541
R15282 iovss.n1105 iovss.n1056 0.00184541
R15283 iovss.n1056 iovss.n961 0.00184541
R15284 iovss.n2752 iovss.n2751 0.00184541
R15285 iovss.n3097 iovss.n1115 0.00184541
R15286 iovss.n3094 iovss.n1115 0.00184541
R15287 iovss.n2900 iovss.n1224 0.00184541
R15288 iovss.n3070 iovss.n2901 0.00184541
R15289 iovss.n2292 iovss.n1731 0.00184541
R15290 iovss.n1803 iovss.n1799 0.00184541
R15291 iovss.n1805 iovss.n1798 0.00184541
R15292 iovss.n1808 iovss.n1797 0.00184541
R15293 iovss.n1810 iovss.n1796 0.00184541
R15294 iovss.n1813 iovss.n1795 0.00184541
R15295 iovss.n1815 iovss.n1794 0.00184541
R15296 iovss.n1818 iovss.n1793 0.00184541
R15297 iovss.n1820 iovss.n1792 0.00184541
R15298 iovss.n1823 iovss.n1791 0.00184541
R15299 iovss.n1827 iovss.n1825 0.00184541
R15300 iovss.n1830 iovss.n1828 0.00184541
R15301 iovss.n1832 iovss.n1831 0.00184541
R15302 iovss.n1835 iovss.n1833 0.00184541
R15303 iovss.n1837 iovss.n1836 0.00184541
R15304 iovss.n1840 iovss.n1838 0.00184541
R15305 iovss.n1843 iovss.n1841 0.00184541
R15306 iovss.n1870 iovss.n1842 0.00184541
R15307 iovss.n1801 iovss.n1800 0.00184541
R15308 iovss.n1807 iovss.n1806 0.00184541
R15309 iovss.n1812 iovss.n1811 0.00184541
R15310 iovss.n1817 iovss.n1816 0.00184541
R15311 iovss.n1822 iovss.n1821 0.00184541
R15312 iovss.n1827 iovss.n1826 0.00184541
R15313 iovss.n1830 iovss.n1829 0.00184541
R15314 iovss.n1835 iovss.n1834 0.00184541
R15315 iovss.n1840 iovss.n1839 0.00184541
R15316 iovss.n1870 iovss.n1869 0.00184541
R15317 iovss.n2095 iovss.n1917 0.00184541
R15318 iovss.n1959 iovss.n1891 0.00184541
R15319 iovss.n2098 iovss.n2096 0.00184541
R15320 iovss.n2101 iovss.n2099 0.00184541
R15321 iovss.n2104 iovss.n2102 0.00184541
R15322 iovss.n2106 iovss.n2105 0.00184541
R15323 iovss.n2109 iovss.n2107 0.00184541
R15324 iovss.n2111 iovss.n2110 0.00184541
R15325 iovss.n2114 iovss.n2112 0.00184541
R15326 iovss.n2116 iovss.n2115 0.00184541
R15327 iovss.n2119 iovss.n2117 0.00184541
R15328 iovss.n2124 iovss.n2122 0.00184541
R15329 iovss.n2129 iovss.n2127 0.00184541
R15330 iovss.n2160 iovss.n2158 0.00184541
R15331 iovss.n2095 iovss.n2094 0.00184541
R15332 iovss.n2098 iovss.n2097 0.00184541
R15333 iovss.n2104 iovss.n2103 0.00184541
R15334 iovss.n2109 iovss.n2108 0.00184541
R15335 iovss.n2114 iovss.n2113 0.00184541
R15336 iovss.n2119 iovss.n2118 0.00184541
R15337 iovss.n2121 iovss.n2120 0.00184541
R15338 iovss.n2124 iovss.n2123 0.00184541
R15339 iovss.n2126 iovss.n2125 0.00184541
R15340 iovss.n2129 iovss.n2128 0.00184541
R15341 iovss.n2131 iovss.n2130 0.00184541
R15342 iovss.n2160 iovss.n2159 0.00184541
R15343 iovss.n2162 iovss.n1944 0.00184541
R15344 iovss.n3079 iovss.n2901 0.00184541
R15345 iovss.n3098 iovss.n3097 0.00184541
R15346 iovss.n3095 iovss.n3094 0.00184541
R15347 iovss.n1105 iovss.n962 0.00184541
R15348 iovss.n3109 iovss.n961 0.00184541
R15349 iovss.n1569 iovss.n1568 0.00184541
R15350 iovss.n1571 iovss.n1570 0.00184541
R15351 iovss.n1573 iovss.n1572 0.00184541
R15352 iovss.n1575 iovss.n1574 0.00184541
R15353 iovss.n1577 iovss.n1576 0.00184541
R15354 iovss.n1579 iovss.n1578 0.00184541
R15355 iovss.n1581 iovss.n1580 0.00184541
R15356 iovss.n1583 iovss.n1582 0.00184541
R15357 iovss.n1585 iovss.n1584 0.00184541
R15358 iovss.n1587 iovss.n1586 0.00184541
R15359 iovss.n1589 iovss.n1588 0.00184541
R15360 iovss.n1591 iovss.n1590 0.00184541
R15361 iovss.n1593 iovss.n1592 0.00184541
R15362 iovss.n1595 iovss.n1594 0.00184541
R15363 iovss.n1598 iovss.n1597 0.00184541
R15364 iovss.n2396 iovss.n1625 0.00184541
R15365 iovss.n2392 iovss.n1571 0.00184541
R15366 iovss.n2391 iovss.n1575 0.00184541
R15367 iovss.n2390 iovss.n1579 0.00184541
R15368 iovss.n2389 iovss.n1583 0.00184541
R15369 iovss.n2388 iovss.n1587 0.00184541
R15370 iovss.n2387 iovss.n1591 0.00184541
R15371 iovss.n2386 iovss.n1593 0.00184541
R15372 iovss.n2385 iovss.n1595 0.00184541
R15373 iovss.n2384 iovss.n1596 0.00184541
R15374 iovss.n2383 iovss.n1598 0.00184541
R15375 iovss.n2382 iovss.n1599 0.00184541
R15376 iovss.n2396 iovss.n1626 0.00184541
R15377 iovss.n2394 iovss.n1550 0.00184541
R15378 iovss.n2886 iovss.n1224 0.00184541
R15379 iovss.n2753 iovss.n2752 0.00184541
R15380 iovss.n767 iovss.n656 0.00184541
R15381 iovss.n767 iovss.n766 0.00184541
R15382 iovss.n730 iovss.n657 0.00184541
R15383 iovss.n728 iovss.n658 0.00184541
R15384 iovss.n725 iovss.n658 0.00184541
R15385 iovss.n726 iovss.n659 0.00184541
R15386 iovss.n723 iovss.n660 0.00184541
R15387 iovss.n720 iovss.n660 0.00184541
R15388 iovss.n721 iovss.n661 0.00184541
R15389 iovss.n718 iovss.n662 0.00184541
R15390 iovss.n715 iovss.n662 0.00184541
R15391 iovss.n716 iovss.n663 0.00184541
R15392 iovss.n713 iovss.n663 0.00184541
R15393 iovss.n3251 iovss.n645 0.00184541
R15394 iovss.n711 iovss.n664 0.00184541
R15395 iovss.n692 iovss.n664 0.00184541
R15396 iovss.n689 iovss.n665 0.00184541
R15397 iovss.n690 iovss.n666 0.00184541
R15398 iovss.n687 iovss.n666 0.00184541
R15399 iovss.n684 iovss.n667 0.00184541
R15400 iovss.n685 iovss.n668 0.00184541
R15401 iovss.n682 iovss.n668 0.00184541
R15402 iovss.n679 iovss.n669 0.00184541
R15403 iovss.n680 iovss.n670 0.00184541
R15404 iovss.n677 iovss.n670 0.00184541
R15405 iovss.n674 iovss.n671 0.00184541
R15406 iovss.n675 iovss.n672 0.00184541
R15407 iovss.n3387 iovss.n286 0.00184541
R15408 iovss.n3387 iovss.n3386 0.00184541
R15409 iovss.n329 iovss.n287 0.00184541
R15410 iovss.n337 iovss.n288 0.00184541
R15411 iovss.n327 iovss.n288 0.00184541
R15412 iovss.n325 iovss.n289 0.00184541
R15413 iovss.n338 iovss.n290 0.00184541
R15414 iovss.n323 iovss.n290 0.00184541
R15415 iovss.n321 iovss.n291 0.00184541
R15416 iovss.n339 iovss.n292 0.00184541
R15417 iovss.n319 iovss.n292 0.00184541
R15418 iovss.n340 iovss.n293 0.00184541
R15419 iovss.n341 iovss.n294 0.00184541
R15420 iovss.n316 iovss.n294 0.00184541
R15421 iovss.n342 iovss.n295 0.00184541
R15422 iovss.n343 iovss.n296 0.00184541
R15423 iovss.n313 iovss.n296 0.00184541
R15424 iovss.n344 iovss.n297 0.00184541
R15425 iovss.n345 iovss.n298 0.00184541
R15426 iovss.n310 iovss.n298 0.00184541
R15427 iovss.n346 iovss.n299 0.00184541
R15428 iovss.n347 iovss.n300 0.00184541
R15429 iovss.n307 iovss.n300 0.00184541
R15430 iovss.n348 iovss.n301 0.00184541
R15431 iovss.n349 iovss.n302 0.00184541
R15432 iovss.n304 iovss.n302 0.00184541
R15433 iovss.n3394 iovss.n265 0.00184541
R15434 iovss.n252 iovss.n203 0.00184541
R15435 iovss.n3416 iovss.n204 0.00184541
R15436 iovss.n249 iovss.n204 0.00184541
R15437 iovss.n3417 iovss.n205 0.00184541
R15438 iovss.n3418 iovss.n206 0.00184541
R15439 iovss.n246 iovss.n206 0.00184541
R15440 iovss.n3419 iovss.n207 0.00184541
R15441 iovss.n244 iovss.n207 0.00184541
R15442 iovss.n3420 iovss.n208 0.00184541
R15443 iovss.n242 iovss.n208 0.00184541
R15444 iovss.n3421 iovss.n209 0.00184541
R15445 iovss.n240 iovss.n209 0.00184541
R15446 iovss.n238 iovss.n210 0.00184541
R15447 iovss.n3429 iovss.n175 0.00184541
R15448 iovss.n3429 iovss.n185 0.00184541
R15449 iovss.n235 iovss.n211 0.00184541
R15450 iovss.n3422 iovss.n212 0.00184541
R15451 iovss.n233 iovss.n212 0.00184541
R15452 iovss.n231 iovss.n213 0.00184541
R15453 iovss.n3423 iovss.n214 0.00184541
R15454 iovss.n229 iovss.n214 0.00184541
R15455 iovss.n227 iovss.n215 0.00184541
R15456 iovss.n3424 iovss.n216 0.00184541
R15457 iovss.n225 iovss.n216 0.00184541
R15458 iovss.n223 iovss.n217 0.00184541
R15459 iovss.n3425 iovss.n218 0.00184541
R15460 iovss.n221 iovss.n218 0.00184541
R15461 iovss.n2716 iovss.n1341 0.00184541
R15462 iovss.n1198 iovss.n912 0.00184541
R15463 iovss.n1310 iovss.n1309 0.00184541
R15464 iovss.n2716 iovss.n1340 0.00184541
R15465 iovss.n2773 iovss.n1310 0.00184541
R15466 iovss.n222 iovss.n221 0.00184541
R15467 iovss.n224 iovss.n223 0.00184541
R15468 iovss.n226 iovss.n225 0.00184541
R15469 iovss.n228 iovss.n227 0.00184541
R15470 iovss.n230 iovss.n229 0.00184541
R15471 iovss.n232 iovss.n231 0.00184541
R15472 iovss.n234 iovss.n233 0.00184541
R15473 iovss.n236 iovss.n235 0.00184541
R15474 iovss.n237 iovss.n185 0.00184541
R15475 iovss.n239 iovss.n238 0.00184541
R15476 iovss.n241 iovss.n240 0.00184541
R15477 iovss.n243 iovss.n242 0.00184541
R15478 iovss.n245 iovss.n244 0.00184541
R15479 iovss.n247 iovss.n246 0.00184541
R15480 iovss.n250 iovss.n249 0.00184541
R15481 iovss.n253 iovss.n252 0.00184541
R15482 iovss.n3425 iovss.n224 0.00184541
R15483 iovss.n3424 iovss.n228 0.00184541
R15484 iovss.n3423 iovss.n232 0.00184541
R15485 iovss.n3422 iovss.n236 0.00184541
R15486 iovss.n239 iovss.n175 0.00184541
R15487 iovss.n3421 iovss.n243 0.00184541
R15488 iovss.n3420 iovss.n245 0.00184541
R15489 iovss.n3419 iovss.n247 0.00184541
R15490 iovss.n3418 iovss.n248 0.00184541
R15491 iovss.n3417 iovss.n250 0.00184541
R15492 iovss.n3416 iovss.n251 0.00184541
R15493 iovss.n305 iovss.n304 0.00184541
R15494 iovss.n308 iovss.n307 0.00184541
R15495 iovss.n311 iovss.n310 0.00184541
R15496 iovss.n314 iovss.n313 0.00184541
R15497 iovss.n317 iovss.n316 0.00184541
R15498 iovss.n320 iovss.n319 0.00184541
R15499 iovss.n322 iovss.n321 0.00184541
R15500 iovss.n324 iovss.n323 0.00184541
R15501 iovss.n326 iovss.n325 0.00184541
R15502 iovss.n328 iovss.n327 0.00184541
R15503 iovss.n330 iovss.n329 0.00184541
R15504 iovss.n3386 iovss.n331 0.00184541
R15505 iovss.n305 iovss.n265 0.00184541
R15506 iovss.n349 iovss.n306 0.00184541
R15507 iovss.n348 iovss.n308 0.00184541
R15508 iovss.n347 iovss.n309 0.00184541
R15509 iovss.n346 iovss.n311 0.00184541
R15510 iovss.n345 iovss.n312 0.00184541
R15511 iovss.n344 iovss.n314 0.00184541
R15512 iovss.n343 iovss.n315 0.00184541
R15513 iovss.n342 iovss.n317 0.00184541
R15514 iovss.n341 iovss.n318 0.00184541
R15515 iovss.n340 iovss.n320 0.00184541
R15516 iovss.n339 iovss.n322 0.00184541
R15517 iovss.n338 iovss.n326 0.00184541
R15518 iovss.n337 iovss.n330 0.00184541
R15519 iovss.n3390 iovss.n286 0.00184541
R15520 iovss.n676 iovss.n674 0.00184541
R15521 iovss.n678 iovss.n677 0.00184541
R15522 iovss.n681 iovss.n679 0.00184541
R15523 iovss.n683 iovss.n682 0.00184541
R15524 iovss.n686 iovss.n684 0.00184541
R15525 iovss.n688 iovss.n687 0.00184541
R15526 iovss.n691 iovss.n689 0.00184541
R15527 iovss.n710 iovss.n692 0.00184541
R15528 iovss.n712 iovss.n645 0.00184541
R15529 iovss.n714 iovss.n713 0.00184541
R15530 iovss.n717 iovss.n715 0.00184541
R15531 iovss.n722 iovss.n720 0.00184541
R15532 iovss.n727 iovss.n725 0.00184541
R15533 iovss.n766 iovss.n731 0.00184541
R15534 iovss.n676 iovss.n675 0.00184541
R15535 iovss.n681 iovss.n680 0.00184541
R15536 iovss.n686 iovss.n685 0.00184541
R15537 iovss.n691 iovss.n690 0.00184541
R15538 iovss.n712 iovss.n711 0.00184541
R15539 iovss.n717 iovss.n716 0.00184541
R15540 iovss.n719 iovss.n718 0.00184541
R15541 iovss.n722 iovss.n721 0.00184541
R15542 iovss.n724 iovss.n723 0.00184541
R15543 iovss.n727 iovss.n726 0.00184541
R15544 iovss.n729 iovss.n728 0.00184541
R15545 iovss.n731 iovss.n730 0.00184541
R15546 iovss.n3246 iovss.n656 0.00184541
R15547 iovss.n3136 iovss.n912 0.00184541
R15548 iovss.n3248 iovss.n742 0.00183951
R15549 iovss.n3334 iovss.n171 0.00182
R15550 iovss.n3321 iovss.n107 0.00182
R15551 iovss.n2211 iovss.n1945 0.00181137
R15552 iovss.n770 iovss.n657 0.00181137
R15553 iovss.n1687 iovss.n1562 0.00177686
R15554 iovss.n856 iovss.n213 0.00177686
R15555 iovss.n2100 iovss.n1958 0.00174235
R15556 iovss.n793 iovss.n669 0.00174235
R15557 iovss.n3134 iovss.n3133 0.00171968
R15558 iovss.n582 iovss.n534 0.00171
R15559 iovss.n2290 iovss.n2288 0.00170784
R15560 iovss.n2273 iovss.n1809 0.00170784
R15561 iovss.n3392 iovss.n333 0.00170784
R15562 iovss.n829 iovss.n309 0.00170784
R15563 iovss.n2180 iovss.n2176 0.0016983
R15564 iovss.n777 iovss.n774 0.0016983
R15565 iovss.n2521 iovss.n1461 0.00167333
R15566 iovss.n2518 iovss.n1465 0.00167333
R15567 iovss.n2240 iovss.n2214 0.00167333
R15568 iovss.n3245 iovss.n742 0.00167333
R15569 iovss.n2564 iovss.n1440 0.0016673
R15570 iovss.n2564 iovss.n1441 0.0016673
R15571 iovss.n2564 iovss.n1448 0.0016673
R15572 iovss.n2564 iovss.n2563 0.0016673
R15573 iovss.n2564 iovss.n1444 0.0016673
R15574 iovss.n2564 iovss.n1443 0.0016673
R15575 iovss.n3253 iovss.n633 0.00165789
R15576 iovss.n3253 iovss.n3252 0.00165789
R15577 iovss.n3363 iovss.n3362 0.00165789
R15578 iovss.n3362 iovss.n3361 0.00165789
R15579 iovss.n3431 iovss.n173 0.00165789
R15580 iovss.n3431 iovss.n3430 0.00165789
R15581 iovss.n2325 iovss.n1564 0.00163882
R15582 iovss.n857 iovss.n215 0.00163882
R15583 iovss.n2244 iovss.n2243 0.00160431
R15584 iovss.n801 iovss.n671 0.00160431
R15585 iovss.n3273 iovss.n432 0.0016
R15586 iovss.n3290 iovss.n446 0.0016
R15587 iovss.n1804 iovss.n1802 0.0015698
R15588 iovss.n830 iovss.n306 0.0015698
R15589 iovss.n3095 iovss.n3083 0.00153529
R15590 iovss.n3136 iovss.n914 0.00153529
R15591 iovss.n2327 iovss.n1566 0.00150078
R15592 iovss.n3070 iovss.n2935 0.00150078
R15593 iovss.n858 iovss.n217 0.00150078
R15594 iovss.n3147 iovss.n886 0.00150078
R15595 iovss.n1112 iovss.n904 0.00149998
R15596 iovss.n1112 iovss.n1111 0.00149998
R15597 iovss.n3102 iovss.n904 0.00149997
R15598 iovss.n3106 iovss.n904 0.00149991
R15599 iovss.n608 iovss.n524 0.00149
R15600 iovss.n1110 iovss.n904 0.0014837
R15601 iovss.n3104 iovss.n3103 0.0014837
R15602 iovss.n1111 iovss.n1110 0.0014837
R15603 iovss.n779 iovss.n778 0.00147778
R15604 iovss.n786 iovss.n779 0.00147778
R15605 iovss.n787 iovss.n786 0.00147778
R15606 iovss.n788 iovss.n787 0.00147778
R15607 iovss.n796 iovss.n788 0.00147778
R15608 iovss.n797 iovss.n796 0.00147778
R15609 iovss.n798 iovss.n797 0.00147778
R15610 iovss.n804 iovss.n798 0.00147778
R15611 iovss.n805 iovss.n804 0.00147778
R15612 iovss.n806 iovss.n805 0.00147778
R15613 iovss.n814 iovss.n806 0.00147778
R15614 iovss.n815 iovss.n814 0.00147778
R15615 iovss.n816 iovss.n815 0.00147778
R15616 iovss.n824 iovss.n816 0.00147778
R15617 iovss.n825 iovss.n824 0.00147778
R15618 iovss.n826 iovss.n825 0.00147778
R15619 iovss.n833 iovss.n826 0.00147778
R15620 iovss.n834 iovss.n833 0.00147778
R15621 iovss.n835 iovss.n834 0.00147778
R15622 iovss.n842 iovss.n835 0.00147778
R15623 iovss.n843 iovss.n842 0.00147778
R15624 iovss.n844 iovss.n843 0.00147778
R15625 iovss.n851 iovss.n844 0.00147778
R15626 iovss.n852 iovss.n851 0.00147778
R15627 iovss.n853 iovss.n852 0.00147778
R15628 iovss.n861 iovss.n853 0.00147778
R15629 iovss.n862 iovss.n861 0.00147778
R15630 iovss.n863 iovss.n862 0.00147778
R15631 iovss.n870 iovss.n863 0.00147778
R15632 iovss.n871 iovss.n870 0.00147778
R15633 iovss.n872 iovss.n871 0.00147778
R15634 iovss.n879 iovss.n872 0.00147778
R15635 iovss.n880 iovss.n879 0.00147778
R15636 iovss.n881 iovss.n880 0.00147778
R15637 iovss.n882 iovss.n881 0.00147778
R15638 iovss.n2184 iovss.n2183 0.00147778
R15639 iovss.n2185 iovss.n2184 0.00147778
R15640 iovss.n2185 iovss.n2173 0.00147778
R15641 iovss.n2192 iovss.n2173 0.00147778
R15642 iovss.n2193 iovss.n2192 0.00147778
R15643 iovss.n2194 iovss.n2193 0.00147778
R15644 iovss.n2196 iovss.n2194 0.00147778
R15645 iovss.n2196 iovss.n2195 0.00147778
R15646 iovss.n2195 iovss.n1888 0.00147778
R15647 iovss.n1888 iovss.n1886 0.00147778
R15648 iovss.n2255 iovss.n1886 0.00147778
R15649 iovss.n2256 iovss.n2255 0.00147778
R15650 iovss.n2257 iovss.n2256 0.00147778
R15651 iovss.n2257 iovss.n1883 0.00147778
R15652 iovss.n2264 iovss.n1883 0.00147778
R15653 iovss.n2265 iovss.n2264 0.00147778
R15654 iovss.n2266 iovss.n2265 0.00147778
R15655 iovss.n2267 iovss.n2266 0.00147778
R15656 iovss.n2267 iovss.n1699 0.00147778
R15657 iovss.n2301 iovss.n1699 0.00147778
R15658 iovss.n2302 iovss.n2301 0.00147778
R15659 iovss.n2303 iovss.n2302 0.00147778
R15660 iovss.n2303 iovss.n1691 0.00147778
R15661 iovss.n2316 iovss.n1691 0.00147778
R15662 iovss.n2317 iovss.n2316 0.00147778
R15663 iovss.n2318 iovss.n2317 0.00147778
R15664 iovss.n2320 iovss.n2318 0.00147778
R15665 iovss.n2320 iovss.n2319 0.00147778
R15666 iovss.n2319 iovss.n1684 0.00147778
R15667 iovss.n2336 iovss.n1684 0.00147778
R15668 iovss.n2337 iovss.n2336 0.00147778
R15669 iovss.n2338 iovss.n2337 0.00147778
R15670 iovss.n2339 iovss.n2338 0.00147778
R15671 iovss.n2340 iovss.n2339 0.00147778
R15672 iovss.n2341 iovss.n2340 0.00147778
R15673 iovss.n2065 iovss.n2026 0.00138
R15674 iovss.n2569 iovss.n1437 0.00138
R15675 iovss.n3330 iovss.n117 0.00138
R15676 iovss.n3323 iovss.n109 0.00138
R15677 iovss.n2355 iovss.n1653 0.00136275
R15678 iovss.n866 iovss.n219 0.00136275
R15679 iovss.n932 iovss.n904 0.00133247
R15680 iovss.n1653 iovss.n1569 0.00132824
R15681 iovss.n866 iovss.n222 0.00132824
R15682 iovss.n567 iovss.n532 0.00127
R15683 iovss.n2293 iovss.n2292 0.00125922
R15684 iovss.n1677 iovss.n962 0.00125922
R15685 iovss.n3394 iovss.n276 0.00125922
R15686 iovss.n949 iovss.n945 0.00125922
R15687 iovss.n46 iovss 0.00125601
R15688 iovss.n47 iovss.n31 0.00120132
R15689 iovss.n2327 iovss.n1573 0.0011902
R15690 iovss.n2935 iovss.n2929 0.0011902
R15691 iovss.n858 iovss.n226 0.0011902
R15692 iovss.n3147 iovss.n3146 0.0011902
R15693 iovss.n3275 iovss.n435 0.00116
R15694 iovss.n3288 iovss.n443 0.00116
R15695 iovss.n1802 iovss.n1798 0.00112118
R15696 iovss.n830 iovss.n301 0.00112118
R15697 iovss.n3138 iovss.n904 0.00109598
R15698 iovss.n2244 iovss.n1891 0.00108667
R15699 iovss.n801 iovss.n678 0.00108667
R15700 iovss.n2325 iovss.n1577 0.00105216
R15701 iovss.n857 iovss.n230 0.00105216
R15702 iovss.n558 iovss.n526 0.00105
R15703 iovss.n2214 iovss.n2162 0.00101765
R15704 iovss.n3246 iovss.n3245 0.00101765
R15705 iovss.n48 iovss.n47 0.00100025
R15706 iovss.n3105 iovss.n3104 0.001
R15707 iovss.n2288 iovss.n1783 0.000983137
R15708 iovss.n2273 iovss.n1796 0.000983137
R15709 iovss.n358 iovss.n333 0.000983137
R15710 iovss.n829 iovss.n299 0.000983137
R15711 iovss.n2101 iovss.n2100 0.000948627
R15712 iovss.n793 iovss.n683 0.000948627
R15713 iovss.n3328 iovss.n115 0.00094
R15714 iovss.n3325 iovss.n111 0.00094
R15715 iovss.n2394 iovss.n1652 0.000914118
R15716 iovss.n1687 iovss.n1581 0.000914118
R15717 iovss.n3427 iovss.n254 0.000914118
R15718 iovss.n856 iovss.n234 0.000914118
R15719 iovss.n48 iovss.n21 0.000902948
R15720 iovss.n48 iovss.n38 0.000888012
R15721 iovss.n48 iovss.n25 0.000888012
R15722 iovss.n2211 iovss.n2131 0.000879608
R15723 iovss.n770 iovss.n729 0.000879608
R15724 iovss.n48 iovss.n37 0.000850673
R15725 iovss.n48 iovss.n24 0.000850673
R15726 iovss.n2285 iovss.n1784 0.000845098
R15727 iovss.n2275 iovss.n1794 0.000845098
R15728 iovss.n809 iovss.n287 0.000845098
R15729 iovss.n821 iovss.n297 0.000845098
R15730 iovss.n593 iovss.n530 0.00083
R15731 iovss.n2201 iovss.n2106 0.000810588
R15732 iovss.n792 iovss.n688 0.000810588
R15733 iovss.n2063 iovss.n2024 0.000793333
R15734 iovss.n2453 iovss.n2452 0.000793333
R15735 iovss.n48 iovss.n22 0.000790931
R15736 iovss.n48 iovss.n35 0.000790931
R15737 iovss.n2296 iovss.n1599 0.000776078
R15738 iovss.n2311 iovss.n1585 0.000776078
R15739 iovss.n838 iovss.n251 0.000776078
R15740 iovss.n848 iovss.n237 0.000776078
R15741 iovss.n2209 iovss.n2126 0.000741569
R15742 iovss.n782 iovss.n724 0.000741569
R15743 iovss.n3277 iovss.n373 0.00072
R15744 iovss.n473 iovss.n440 0.00072
R15745 iovss.n48 iovss.n44 0.000708786
R15746 iovss.n2283 iovss.n1786 0.000707059
R15747 iovss.n2277 iovss.n1792 0.000707059
R15748 iovss.n810 iovss.n289 0.000707059
R15749 iovss.n820 iovss.n295 0.000707059
R15750 iovss.n49 iovss.n48 0.000676426
R15751 iovss.n2203 iovss.n2111 0.000672549
R15752 iovss.n3080 iovss.n2900 0.000672549
R15753 iovss.n791 iovss.n710 0.000672549
R15754 iovss.n1312 iovss.n885 0.000672549
R15755 iovss.n1695 iovss.n1596 0.000638039
R15756 iovss.n2309 iovss.n1589 0.000638039
R15757 iovss.n839 iovss.n248 0.000638039
R15758 iovss.n847 iovss.n241 0.000638039
R15759 iovss.n595 iovss.n528 0.00061
R15760 iovss.n2207 iovss.n2121 0.000603529
R15761 iovss.n783 iovss.n719 0.000603529
R15762 iovss.n46 iovss 0.000570408
R15763 iovss.n2281 iovss.n1788 0.00056902
R15764 iovss.n2279 iovss.n1790 0.00056902
R15765 iovss.n811 iovss.n291 0.00056902
R15766 iovss.n819 iovss.n293 0.00056902
R15767 iovss.n48 iovss.n23 0.000564409
R15768 iovss.n48 iovss.n36 0.000564409
R15769 iovss.n2205 iovss.n2116 0.00053451
R15770 iovss.n714 iovss.n635 0.00053451
R15771 iovdd.n1307 iovdd.n43 17.0005
R15772 iovdd.n1307 iovdd.n5 17.0005
R15773 iovdd.n49 iovdd.n43 17.0005
R15774 iovdd.n49 iovdd.n4 17.0005
R15775 iovdd.n1359 iovdd.n49 17.0005
R15776 iovdd.n49 iovdd.n42 17.0005
R15777 iovdd.n49 iovdd.n40 17.0005
R15778 iovdd.n49 iovdd.n39 17.0005
R15779 iovdd.n49 iovdd.n37 17.0005
R15780 iovdd.n49 iovdd.n36 17.0005
R15781 iovdd.n49 iovdd.n34 17.0005
R15782 iovdd.n49 iovdd.n33 17.0005
R15783 iovdd.n49 iovdd.n31 17.0005
R15784 iovdd.n49 iovdd.n30 17.0005
R15785 iovdd.n49 iovdd.n28 17.0005
R15786 iovdd.n49 iovdd.n27 17.0005
R15787 iovdd.n49 iovdd.n23 17.0005
R15788 iovdd.n49 iovdd.n22 17.0005
R15789 iovdd.n49 iovdd.n20 17.0005
R15790 iovdd.n49 iovdd.n19 17.0005
R15791 iovdd.n49 iovdd.n17 17.0005
R15792 iovdd.n49 iovdd.n16 17.0005
R15793 iovdd.n49 iovdd.n13 17.0005
R15794 iovdd.n49 iovdd.n12 17.0005
R15795 iovdd.n49 iovdd.n11 17.0005
R15796 iovdd.n49 iovdd.n10 17.0005
R15797 iovdd.n49 iovdd.n9 17.0005
R15798 iovdd.n1229 iovdd.n49 17.0005
R15799 iovdd.n49 iovdd.n7 17.0005
R15800 iovdd.n49 iovdd.n5 17.0005
R15801 iovdd.n1313 iovdd.n272 9.0005
R15802 iovdd.n1313 iovdd.n273 9.0005
R15803 iovdd.n547 iovdd.n479 9.0005
R15804 iovdd.n547 iovdd.n483 9.0005
R15805 iovdd.n547 iovdd.n476 9.0005
R15806 iovdd.n547 iovdd.n486 9.0005
R15807 iovdd.n547 iovdd.n474 9.0005
R15808 iovdd.n547 iovdd.n489 9.0005
R15809 iovdd.n547 iovdd.n472 9.0005
R15810 iovdd.n547 iovdd.n492 9.0005
R15811 iovdd.n547 iovdd.n470 9.0005
R15812 iovdd.n547 iovdd.n495 9.0005
R15813 iovdd.n547 iovdd.n468 9.0005
R15814 iovdd.n547 iovdd.n498 9.0005
R15815 iovdd.n547 iovdd.n466 9.0005
R15816 iovdd.n547 iovdd.n501 9.0005
R15817 iovdd.n547 iovdd.n464 9.0005
R15818 iovdd.n547 iovdd.n504 9.0005
R15819 iovdd.n547 iovdd.n462 9.0005
R15820 iovdd.n547 iovdd.n507 9.0005
R15821 iovdd.n547 iovdd.n460 9.0005
R15822 iovdd.n547 iovdd.n510 9.0005
R15823 iovdd.n547 iovdd.n458 9.0005
R15824 iovdd.n547 iovdd.n513 9.0005
R15825 iovdd.n547 iovdd.n456 9.0005
R15826 iovdd.n547 iovdd.n516 9.0005
R15827 iovdd.n547 iovdd.n454 9.0005
R15828 iovdd.n547 iovdd.n519 9.0005
R15829 iovdd.n547 iovdd.n452 9.0005
R15830 iovdd.n547 iovdd.n522 9.0005
R15831 iovdd.n547 iovdd.n450 9.0005
R15832 iovdd.n547 iovdd.n525 9.0005
R15833 iovdd.n547 iovdd.n448 9.0005
R15834 iovdd.n547 iovdd.n528 9.0005
R15835 iovdd.n547 iovdd.n446 9.0005
R15836 iovdd.n547 iovdd.n531 9.0005
R15837 iovdd.n547 iovdd.n444 9.0005
R15838 iovdd.n547 iovdd.n534 9.0005
R15839 iovdd.n547 iovdd.n442 9.0005
R15840 iovdd.n547 iovdd.n537 9.0005
R15841 iovdd.n547 iovdd.n440 9.0005
R15842 iovdd.n547 iovdd.n540 9.0005
R15843 iovdd.n547 iovdd.n438 9.0005
R15844 iovdd.n547 iovdd.n543 9.0005
R15845 iovdd.n547 iovdd.n436 9.0005
R15846 iovdd.n547 iovdd.n546 9.0005
R15847 iovdd.n547 iovdd.n434 9.0005
R15848 iovdd.n1313 iovdd.n1312 9.0005
R15849 iovdd.n1223 iovdd.n862 9.0005
R15850 iovdd.n1221 iovdd.n862 9.0005
R15851 iovdd.n1218 iovdd.n862 9.0005
R15852 iovdd.n1221 iovdd.n1136 9.0005
R15853 iovdd.n1221 iovdd.n1138 9.0005
R15854 iovdd.n1221 iovdd.n1134 9.0005
R15855 iovdd.n1221 iovdd.n1140 9.0005
R15856 iovdd.n1221 iovdd.n1132 9.0005
R15857 iovdd.n1221 iovdd.n1142 9.0005
R15858 iovdd.n1221 iovdd.n1130 9.0005
R15859 iovdd.n1221 iovdd.n1144 9.0005
R15860 iovdd.n1221 iovdd.n1128 9.0005
R15861 iovdd.n1221 iovdd.n1146 9.0005
R15862 iovdd.n1221 iovdd.n1126 9.0005
R15863 iovdd.n1221 iovdd.n1148 9.0005
R15864 iovdd.n1221 iovdd.n1124 9.0005
R15865 iovdd.n1221 iovdd.n1150 9.0005
R15866 iovdd.n1221 iovdd.n1122 9.0005
R15867 iovdd.n1221 iovdd.n1152 9.0005
R15868 iovdd.n1221 iovdd.n1120 9.0005
R15869 iovdd.n1221 iovdd.n1154 9.0005
R15870 iovdd.n1221 iovdd.n1118 9.0005
R15871 iovdd.n1221 iovdd.n1156 9.0005
R15872 iovdd.n1221 iovdd.n1116 9.0005
R15873 iovdd.n1221 iovdd.n1158 9.0005
R15874 iovdd.n1221 iovdd.n1114 9.0005
R15875 iovdd.n1221 iovdd.n1160 9.0005
R15876 iovdd.n1221 iovdd.n1112 9.0005
R15877 iovdd.n1221 iovdd.n1162 9.0005
R15878 iovdd.n1221 iovdd.n1110 9.0005
R15879 iovdd.n1221 iovdd.n1164 9.0005
R15880 iovdd.n1221 iovdd.n1108 9.0005
R15881 iovdd.n1221 iovdd.n1166 9.0005
R15882 iovdd.n1221 iovdd.n1106 9.0005
R15883 iovdd.n1221 iovdd.n1168 9.0005
R15884 iovdd.n1221 iovdd.n1104 9.0005
R15885 iovdd.n1221 iovdd.n1170 9.0005
R15886 iovdd.n1221 iovdd.n1102 9.0005
R15887 iovdd.n1221 iovdd.n1172 9.0005
R15888 iovdd.n1221 iovdd.n1100 9.0005
R15889 iovdd.n1221 iovdd.n1174 9.0005
R15890 iovdd.n1221 iovdd.n1098 9.0005
R15891 iovdd.n1221 iovdd.n1176 9.0005
R15892 iovdd.n1221 iovdd.n1096 9.0005
R15893 iovdd.n1221 iovdd.n1178 9.0005
R15894 iovdd.n1221 iovdd.n1094 9.0005
R15895 iovdd.n1221 iovdd.n1180 9.0005
R15896 iovdd.n1221 iovdd.n1092 9.0005
R15897 iovdd.n1221 iovdd.n1220 9.0005
R15898 iovdd.n1220 iovdd.n1218 9.0005
R15899 iovdd.n1218 iovdd.n860 9.0005
R15900 iovdd.n1221 iovdd.n860 9.0005
R15901 iovdd.n297 iovdd.n290 9.0005
R15902 iovdd.n297 iovdd.n275 9.0005
R15903 iovdd.n1311 iovdd.n297 9.0005
R15904 iovdd.n1225 iovdd.n860 9.0005
R15905 iovdd.n1227 iovdd.n860 9.0005
R15906 iovdd.n863 iovdd.n860 9.0005
R15907 iovdd.n1312 iovdd.n290 9.0005
R15908 iovdd.n1312 iovdd.n275 9.0005
R15909 iovdd.n1312 iovdd.n1311 9.0005
R15910 iovdd.n1226 iovdd.n1225 9.0005
R15911 iovdd.n1226 iovdd.n863 9.0005
R15912 iovdd.n1227 iovdd.n1226 9.0005
R15913 iovdd.n1357 iovdd.n113 9.0005
R15914 iovdd.n113 iovdd.n111 9.0005
R15915 iovdd.n1357 iovdd.n1356 9.0005
R15916 iovdd.n1355 iovdd.n165 9.0005
R15917 iovdd.n1355 iovdd.n168 9.0005
R15918 iovdd.n1355 iovdd.n164 9.0005
R15919 iovdd.n1355 iovdd.n171 9.0005
R15920 iovdd.n1355 iovdd.n162 9.0005
R15921 iovdd.n1355 iovdd.n174 9.0005
R15922 iovdd.n1355 iovdd.n160 9.0005
R15923 iovdd.n1355 iovdd.n177 9.0005
R15924 iovdd.n1355 iovdd.n158 9.0005
R15925 iovdd.n1355 iovdd.n180 9.0005
R15926 iovdd.n1355 iovdd.n156 9.0005
R15927 iovdd.n1355 iovdd.n183 9.0005
R15928 iovdd.n1355 iovdd.n154 9.0005
R15929 iovdd.n1355 iovdd.n186 9.0005
R15930 iovdd.n1355 iovdd.n152 9.0005
R15931 iovdd.n1355 iovdd.n189 9.0005
R15932 iovdd.n1355 iovdd.n150 9.0005
R15933 iovdd.n1355 iovdd.n192 9.0005
R15934 iovdd.n1355 iovdd.n148 9.0005
R15935 iovdd.n1355 iovdd.n195 9.0005
R15936 iovdd.n1355 iovdd.n146 9.0005
R15937 iovdd.n1355 iovdd.n198 9.0005
R15938 iovdd.n1355 iovdd.n144 9.0005
R15939 iovdd.n1355 iovdd.n201 9.0005
R15940 iovdd.n1355 iovdd.n142 9.0005
R15941 iovdd.n1355 iovdd.n204 9.0005
R15942 iovdd.n1355 iovdd.n140 9.0005
R15943 iovdd.n1355 iovdd.n207 9.0005
R15944 iovdd.n1355 iovdd.n138 9.0005
R15945 iovdd.n1355 iovdd.n210 9.0005
R15946 iovdd.n1355 iovdd.n136 9.0005
R15947 iovdd.n1355 iovdd.n213 9.0005
R15948 iovdd.n1355 iovdd.n134 9.0005
R15949 iovdd.n1355 iovdd.n216 9.0005
R15950 iovdd.n1355 iovdd.n132 9.0005
R15951 iovdd.n1355 iovdd.n219 9.0005
R15952 iovdd.n1355 iovdd.n130 9.0005
R15953 iovdd.n1355 iovdd.n222 9.0005
R15954 iovdd.n1355 iovdd.n128 9.0005
R15955 iovdd.n1355 iovdd.n225 9.0005
R15956 iovdd.n1355 iovdd.n126 9.0005
R15957 iovdd.n1355 iovdd.n228 9.0005
R15958 iovdd.n1355 iovdd.n124 9.0005
R15959 iovdd.n1355 iovdd.n231 9.0005
R15960 iovdd.n1355 iovdd.n122 9.0005
R15961 iovdd.n1355 iovdd.n234 9.0005
R15962 iovdd.n1355 iovdd.n120 9.0005
R15963 iovdd.n1354 iovdd.n1353 9.0005
R15964 iovdd.n1355 iovdd.n1354 9.0005
R15965 iovdd.n1356 iovdd.n115 9.0005
R15966 iovdd.n1356 iovdd.n1355 9.0005
R15967 iovdd.n1355 iovdd.n113 9.0005
R15968 iovdd.n1356 iovdd.n111 9.0005
R15969 iovdd.n1301 iovdd.n1300 9.0005
R15970 iovdd.n1304 iovdd.n400 9.0005
R15971 iovdd.n1304 iovdd.n404 9.0005
R15972 iovdd.n1304 iovdd.n398 9.0005
R15973 iovdd.n1304 iovdd.n407 9.0005
R15974 iovdd.n1304 iovdd.n396 9.0005
R15975 iovdd.n1304 iovdd.n410 9.0005
R15976 iovdd.n1304 iovdd.n394 9.0005
R15977 iovdd.n1304 iovdd.n1303 9.0005
R15978 iovdd.n1304 iovdd.n392 9.0005
R15979 iovdd.n1305 iovdd.n389 9.0005
R15980 iovdd.n1305 iovdd.n1304 9.0005
R15981 iovdd.n1264 iovdd.n424 9.0005
R15982 iovdd.n1261 iovdd.n424 9.0005
R15983 iovdd.n1261 iovdd.n1251 9.0005
R15984 iovdd.n1261 iovdd.n1248 9.0005
R15985 iovdd.n1261 iovdd.n1254 9.0005
R15986 iovdd.n1261 iovdd.n1246 9.0005
R15987 iovdd.n1261 iovdd.n1257 9.0005
R15988 iovdd.n1261 iovdd.n1244 9.0005
R15989 iovdd.n1261 iovdd.n1260 9.0005
R15990 iovdd.n1261 iovdd.n1242 9.0005
R15991 iovdd.n1262 iovdd.n1261 9.0005
R15992 iovdd.n1261 iovdd.n565 9.0005
R15993 iovdd.n1264 iovdd.n388 9.0005
R15994 iovdd.n1261 iovdd.n388 9.0005
R15995 iovdd.n1236 iovdd.n771 9.0005
R15996 iovdd.n1233 iovdd.n771 9.0005
R15997 iovdd.n1233 iovdd.n786 9.0005
R15998 iovdd.n1233 iovdd.n784 9.0005
R15999 iovdd.n1233 iovdd.n788 9.0005
R16000 iovdd.n1233 iovdd.n783 9.0005
R16001 iovdd.n1233 iovdd.n1232 9.0005
R16002 iovdd.n1233 iovdd.n782 9.0005
R16003 iovdd.n1234 iovdd.n1233 9.0005
R16004 iovdd.n1233 iovdd.n778 9.0005
R16005 iovdd.n1237 iovdd.n1236 9.0005
R16006 iovdd.n774 iovdd.n773 9.0005
R16007 iovdd.n1307 iovdd.n47 8.501
R16008 iovdd.n1307 iovdd.n386 8.501
R16009 iovdd.n1307 iovdd.n385 8.501
R16010 iovdd.n1307 iovdd.n384 8.501
R16011 iovdd.n1307 iovdd.n383 8.501
R16012 iovdd.n1307 iovdd.n382 8.501
R16013 iovdd.n1307 iovdd.n362 8.501
R16014 iovdd.n1308 iovdd.n1307 8.501
R16015 iovdd.n1307 iovdd.n381 8.501
R16016 iovdd.n1307 iovdd.n380 8.501
R16017 iovdd.n1307 iovdd.n379 8.501
R16018 iovdd.n1307 iovdd.n378 8.501
R16019 iovdd.n1307 iovdd.n377 8.501
R16020 iovdd.n1307 iovdd.n376 8.501
R16021 iovdd.n375 iovdd.n374 8.501
R16022 iovdd.n375 iovdd.n48 8.501
R16023 iovdd.n375 iovdd.n373 8.501
R16024 iovdd.n375 iovdd.n372 8.501
R16025 iovdd.n375 iovdd.n371 8.501
R16026 iovdd.n375 iovdd.n370 8.501
R16027 iovdd.n375 iovdd.n369 8.501
R16028 iovdd.n375 iovdd.n368 8.501
R16029 iovdd.n375 iovdd.n367 8.501
R16030 iovdd.n375 iovdd.n366 8.501
R16031 iovdd.n375 iovdd.n365 8.501
R16032 iovdd.n375 iovdd.n364 8.501
R16033 iovdd.n857 iovdd.n375 8.501
R16034 iovdd.n375 iovdd.n363 8.501
R16035 iovdd.n1309 iovdd.n375 8.5005
R16036 iovdd.n1309 iovdd.n49 8.5005
R16037 iovdd.n1360 iovdd.n44 5.66866
R16038 iovdd.n858 iovdd.n6 5.66767
R16039 iovdd.n1309 iovdd.n359 5.66717
R16040 iovdd.n1309 iovdd.n357 5.66717
R16041 iovdd.n1309 iovdd.n356 5.66717
R16042 iovdd.n1309 iovdd.n354 5.66717
R16043 iovdd.n1309 iovdd.n352 5.66717
R16044 iovdd.n1309 iovdd.n350 5.66717
R16045 iovdd.n1309 iovdd.n348 5.66717
R16046 iovdd.n1309 iovdd.n347 5.66717
R16047 iovdd.n1309 iovdd.n345 5.66717
R16048 iovdd.n1309 iovdd.n343 5.66717
R16049 iovdd.n1309 iovdd.n341 5.66717
R16050 iovdd.n1309 iovdd.n339 5.66717
R16051 iovdd.n1309 iovdd.n338 5.66717
R16052 iovdd.n1309 iovdd.n336 5.66717
R16053 iovdd.n1309 iovdd.n334 5.66717
R16054 iovdd.n1309 iovdd.n332 5.66717
R16055 iovdd.n1309 iovdd.n330 5.66717
R16056 iovdd.n1309 iovdd.n329 5.66717
R16057 iovdd.n1309 iovdd.n327 5.66717
R16058 iovdd.n1309 iovdd.n325 5.66717
R16059 iovdd.n1309 iovdd.n323 5.66717
R16060 iovdd.n1309 iovdd.n322 5.66717
R16061 iovdd.n1309 iovdd.n320 5.66717
R16062 iovdd.n1309 iovdd.n318 5.66717
R16063 iovdd.n1309 iovdd.n316 5.66717
R16064 iovdd.n1309 iovdd.n314 5.66717
R16065 iovdd.n1309 iovdd.n313 5.66717
R16066 iovdd.n1309 iovdd.n311 5.66717
R16067 iovdd.n1309 iovdd.n309 5.66717
R16068 iovdd.n1309 iovdd.n307 5.66717
R16069 iovdd.n1309 iovdd.n305 5.66717
R16070 iovdd.n1309 iovdd.n304 5.66717
R16071 iovdd.n1309 iovdd.n302 5.66717
R16072 iovdd.n1309 iovdd.n299 5.66717
R16073 iovdd.n1309 iovdd.n361 5.66717
R16074 iovdd.n1229 iovdd.n567 5.66717
R16075 iovdd.n1229 iovdd.n854 5.66717
R16076 iovdd.n1230 iovdd.n1229 5.66717
R16077 iovdd.n1229 iovdd.n852 5.66717
R16078 iovdd.n1229 iovdd.n848 5.66717
R16079 iovdd.n1229 iovdd.n844 5.66717
R16080 iovdd.n1229 iovdd.n842 5.66717
R16081 iovdd.n1229 iovdd.n840 5.66717
R16082 iovdd.n1229 iovdd.n839 5.66717
R16083 iovdd.n1229 iovdd.n837 5.66717
R16084 iovdd.n1229 iovdd.n835 5.66717
R16085 iovdd.n1229 iovdd.n833 5.66717
R16086 iovdd.n1229 iovdd.n831 5.66717
R16087 iovdd.n1229 iovdd.n830 5.66717
R16088 iovdd.n1229 iovdd.n828 5.66717
R16089 iovdd.n1229 iovdd.n826 5.66717
R16090 iovdd.n1229 iovdd.n824 5.66717
R16091 iovdd.n1229 iovdd.n823 5.66717
R16092 iovdd.n1229 iovdd.n821 5.66717
R16093 iovdd.n1229 iovdd.n819 5.66717
R16094 iovdd.n1229 iovdd.n817 5.66717
R16095 iovdd.n1229 iovdd.n815 5.66717
R16096 iovdd.n1229 iovdd.n814 5.66717
R16097 iovdd.n1229 iovdd.n812 5.66717
R16098 iovdd.n1229 iovdd.n810 5.66717
R16099 iovdd.n1229 iovdd.n808 5.66717
R16100 iovdd.n1229 iovdd.n806 5.66717
R16101 iovdd.n1229 iovdd.n805 5.66717
R16102 iovdd.n1229 iovdd.n803 5.66717
R16103 iovdd.n1229 iovdd.n801 5.66717
R16104 iovdd.n1229 iovdd.n799 5.66717
R16105 iovdd.n1229 iovdd.n797 5.66717
R16106 iovdd.n1229 iovdd.n796 5.66717
R16107 iovdd.n1229 iovdd.n794 5.66717
R16108 iovdd.n1229 iovdd.n792 5.66717
R16109 iovdd.t0 iovdd.n43 5.66717
R16110 iovdd.t0 iovdd.n4 5.66717
R16111 iovdd.t0 iovdd.n42 5.66717
R16112 iovdd.t0 iovdd.n40 5.66717
R16113 iovdd.t0 iovdd.n39 5.66717
R16114 iovdd.t0 iovdd.n37 5.66717
R16115 iovdd.t0 iovdd.n36 5.66717
R16116 iovdd.t0 iovdd.n34 5.66717
R16117 iovdd.t0 iovdd.n33 5.66717
R16118 iovdd.t0 iovdd.n31 5.66717
R16119 iovdd.t0 iovdd.n30 5.66717
R16120 iovdd.t0 iovdd.n28 5.66717
R16121 iovdd.t0 iovdd.n27 5.66717
R16122 iovdd.t0 iovdd.n23 5.66717
R16123 iovdd.t0 iovdd.n22 5.66717
R16124 iovdd.t0 iovdd.n20 5.66717
R16125 iovdd.t0 iovdd.n19 5.66717
R16126 iovdd.t0 iovdd.n17 5.66717
R16127 iovdd.t0 iovdd.n16 5.66717
R16128 iovdd.t0 iovdd.n13 5.66717
R16129 iovdd.t0 iovdd.n12 5.66717
R16130 iovdd.t0 iovdd.n11 5.66717
R16131 iovdd.t0 iovdd.n10 5.66717
R16132 iovdd.t0 iovdd.n9 5.66717
R16133 iovdd.t0 iovdd.n7 5.66717
R16134 iovdd.t0 iovdd.n5 5.66717
R16135 iovdd.n1359 iovdd.n108 5.66717
R16136 iovdd.n1359 iovdd.n106 5.66717
R16137 iovdd.n1359 iovdd.n105 5.66717
R16138 iovdd.n1359 iovdd.n103 5.66717
R16139 iovdd.n1359 iovdd.n101 5.66717
R16140 iovdd.n1359 iovdd.n99 5.66717
R16141 iovdd.n1359 iovdd.n97 5.66717
R16142 iovdd.n1359 iovdd.n96 5.66717
R16143 iovdd.n1359 iovdd.n94 5.66717
R16144 iovdd.n1359 iovdd.n92 5.66717
R16145 iovdd.n1359 iovdd.n90 5.66717
R16146 iovdd.n1359 iovdd.n88 5.66717
R16147 iovdd.n1359 iovdd.n87 5.66717
R16148 iovdd.n1359 iovdd.n85 5.66717
R16149 iovdd.n1359 iovdd.n83 5.66717
R16150 iovdd.n1359 iovdd.n81 5.66717
R16151 iovdd.n1359 iovdd.n80 5.66717
R16152 iovdd.n1359 iovdd.n78 5.66717
R16153 iovdd.n1359 iovdd.n76 5.66717
R16154 iovdd.n1359 iovdd.n74 5.66717
R16155 iovdd.n1359 iovdd.n72 5.66717
R16156 iovdd.n1359 iovdd.n71 5.66717
R16157 iovdd.n1359 iovdd.n69 5.66717
R16158 iovdd.n1359 iovdd.n67 5.66717
R16159 iovdd.n1359 iovdd.n65 5.66717
R16160 iovdd.n1359 iovdd.n63 5.66717
R16161 iovdd.n1359 iovdd.n62 5.66717
R16162 iovdd.n1359 iovdd.n60 5.66717
R16163 iovdd.n1359 iovdd.n58 5.66717
R16164 iovdd.n1359 iovdd.n56 5.66717
R16165 iovdd.n1359 iovdd.n54 5.66717
R16166 iovdd.n1359 iovdd.n53 5.66717
R16167 iovdd.n1359 iovdd.n51 5.66717
R16168 iovdd.n1359 iovdd.n46 5.66717
R16169 iovdd.n1359 iovdd.n110 5.66717
R16170 iovdd.n1359 iovdd.n45 5.66717
R16171 iovdd.n1359 iovdd.n1358 5.66717
R16172 iovdd.n289 iovdd.n288 5.66717
R16173 iovdd.n288 iovdd.n277 5.66717
R16174 iovdd.n1310 iovdd.n1309 5.66717
R16175 iovdd.n3 iovdd.n0 5.66717
R16176 iovdd.n861 iovdd.n3 5.66717
R16177 iovdd.n1229 iovdd.n1228 5.66717
R16178 iovdd.n550 iovdd.n548 4.50058
R16179 iovdd.n297 iovdd.n248 4.50058
R16180 iovdd.n1222 iovdd.n1089 4.50058
R16181 iovdd.n1226 iovdd.n864 4.50058
R16182 iovdd.n1329 iovdd.n113 4.50058
R16183 iovdd.n1297 iovdd.n1296 4.50058
R16184 iovdd.n781 iovdd.n387 4.50058
R16185 iovdd.n547 iovdd.n480 4.49246
R16186 iovdd.n477 iovdd.n431 4.49246
R16187 iovdd.n1313 iovdd.n271 4.49246
R16188 iovdd.n481 iovdd.n431 4.49246
R16189 iovdd.n1313 iovdd.n270 4.49246
R16190 iovdd.n484 iovdd.n431 4.49246
R16191 iovdd.n1313 iovdd.n269 4.49246
R16192 iovdd.n487 iovdd.n431 4.49246
R16193 iovdd.n1313 iovdd.n268 4.49246
R16194 iovdd.n490 iovdd.n431 4.49246
R16195 iovdd.n1313 iovdd.n267 4.49246
R16196 iovdd.n493 iovdd.n431 4.49246
R16197 iovdd.n1313 iovdd.n266 4.49246
R16198 iovdd.n496 iovdd.n431 4.49246
R16199 iovdd.n1313 iovdd.n265 4.49246
R16200 iovdd.n499 iovdd.n431 4.49246
R16201 iovdd.n1313 iovdd.n264 4.49246
R16202 iovdd.n502 iovdd.n431 4.49246
R16203 iovdd.n1313 iovdd.n263 4.49246
R16204 iovdd.n505 iovdd.n431 4.49246
R16205 iovdd.n1313 iovdd.n262 4.49246
R16206 iovdd.n508 iovdd.n431 4.49246
R16207 iovdd.n1313 iovdd.n261 4.49246
R16208 iovdd.n511 iovdd.n431 4.49246
R16209 iovdd.n1313 iovdd.n260 4.49246
R16210 iovdd.n514 iovdd.n431 4.49246
R16211 iovdd.n1313 iovdd.n259 4.49246
R16212 iovdd.n517 iovdd.n431 4.49246
R16213 iovdd.n1313 iovdd.n258 4.49246
R16214 iovdd.n520 iovdd.n431 4.49246
R16215 iovdd.n1313 iovdd.n257 4.49246
R16216 iovdd.n523 iovdd.n431 4.49246
R16217 iovdd.n1313 iovdd.n256 4.49246
R16218 iovdd.n526 iovdd.n431 4.49246
R16219 iovdd.n1313 iovdd.n255 4.49246
R16220 iovdd.n529 iovdd.n431 4.49246
R16221 iovdd.n1313 iovdd.n254 4.49246
R16222 iovdd.n532 iovdd.n431 4.49246
R16223 iovdd.n1313 iovdd.n253 4.49246
R16224 iovdd.n535 iovdd.n431 4.49246
R16225 iovdd.n1313 iovdd.n252 4.49246
R16226 iovdd.n538 iovdd.n431 4.49246
R16227 iovdd.n1313 iovdd.n251 4.49246
R16228 iovdd.n541 iovdd.n431 4.49246
R16229 iovdd.n1313 iovdd.n250 4.49246
R16230 iovdd.n544 iovdd.n431 4.49246
R16231 iovdd.n1313 iovdd.n249 4.49246
R16232 iovdd.n431 iovdd.n274 4.49246
R16233 iovdd.n547 iovdd.n276 4.49246
R16234 iovdd.n1218 iovdd.n1217 4.49246
R16235 iovdd.n1223 iovdd.n1087 4.49246
R16236 iovdd.n1218 iovdd.n1216 4.49246
R16237 iovdd.n1223 iovdd.n1086 4.49246
R16238 iovdd.n1218 iovdd.n1215 4.49246
R16239 iovdd.n1223 iovdd.n1085 4.49246
R16240 iovdd.n1218 iovdd.n1214 4.49246
R16241 iovdd.n1223 iovdd.n1084 4.49246
R16242 iovdd.n1218 iovdd.n1213 4.49246
R16243 iovdd.n1223 iovdd.n1083 4.49246
R16244 iovdd.n1218 iovdd.n1212 4.49246
R16245 iovdd.n1223 iovdd.n1082 4.49246
R16246 iovdd.n1218 iovdd.n1211 4.49246
R16247 iovdd.n1223 iovdd.n1081 4.49246
R16248 iovdd.n1218 iovdd.n1210 4.49246
R16249 iovdd.n1223 iovdd.n1080 4.49246
R16250 iovdd.n1218 iovdd.n1209 4.49246
R16251 iovdd.n1223 iovdd.n1079 4.49246
R16252 iovdd.n1218 iovdd.n1208 4.49246
R16253 iovdd.n1223 iovdd.n1078 4.49246
R16254 iovdd.n1218 iovdd.n1207 4.49246
R16255 iovdd.n1223 iovdd.n1077 4.49246
R16256 iovdd.n1218 iovdd.n1206 4.49246
R16257 iovdd.n1223 iovdd.n1076 4.49246
R16258 iovdd.n1218 iovdd.n1205 4.49246
R16259 iovdd.n1223 iovdd.n1075 4.49246
R16260 iovdd.n1218 iovdd.n1204 4.49246
R16261 iovdd.n1223 iovdd.n1074 4.49246
R16262 iovdd.n1218 iovdd.n1203 4.49246
R16263 iovdd.n1223 iovdd.n1073 4.49246
R16264 iovdd.n1218 iovdd.n1202 4.49246
R16265 iovdd.n1223 iovdd.n1072 4.49246
R16266 iovdd.n1218 iovdd.n1201 4.49246
R16267 iovdd.n1223 iovdd.n1071 4.49246
R16268 iovdd.n1218 iovdd.n1200 4.49246
R16269 iovdd.n1223 iovdd.n1070 4.49246
R16270 iovdd.n1218 iovdd.n1199 4.49246
R16271 iovdd.n1223 iovdd.n1069 4.49246
R16272 iovdd.n1218 iovdd.n1198 4.49246
R16273 iovdd.n1223 iovdd.n1068 4.49246
R16274 iovdd.n1218 iovdd.n1197 4.49246
R16275 iovdd.n1223 iovdd.n1067 4.49246
R16276 iovdd.n1218 iovdd.n1196 4.49246
R16277 iovdd.n1223 iovdd.n1066 4.49246
R16278 iovdd.n1218 iovdd.n1195 4.49246
R16279 iovdd.n1223 iovdd.n1065 4.49246
R16280 iovdd.n1224 iovdd.n1223 4.49246
R16281 iovdd.n117 iovdd.n116 4.49246
R16282 iovdd.n1353 iovdd.n114 4.49246
R16283 iovdd.n166 iovdd.n115 4.49246
R16284 iovdd.n1353 iovdd.n1330 4.49246
R16285 iovdd.n169 iovdd.n115 4.49246
R16286 iovdd.n1353 iovdd.n1331 4.49246
R16287 iovdd.n172 iovdd.n115 4.49246
R16288 iovdd.n1353 iovdd.n1332 4.49246
R16289 iovdd.n175 iovdd.n115 4.49246
R16290 iovdd.n1353 iovdd.n1333 4.49246
R16291 iovdd.n178 iovdd.n115 4.49246
R16292 iovdd.n1353 iovdd.n1334 4.49246
R16293 iovdd.n181 iovdd.n115 4.49246
R16294 iovdd.n1353 iovdd.n1335 4.49246
R16295 iovdd.n184 iovdd.n115 4.49246
R16296 iovdd.n1353 iovdd.n1336 4.49246
R16297 iovdd.n187 iovdd.n115 4.49246
R16298 iovdd.n1353 iovdd.n1337 4.49246
R16299 iovdd.n190 iovdd.n115 4.49246
R16300 iovdd.n1353 iovdd.n1338 4.49246
R16301 iovdd.n193 iovdd.n115 4.49246
R16302 iovdd.n1353 iovdd.n1339 4.49246
R16303 iovdd.n196 iovdd.n115 4.49246
R16304 iovdd.n1353 iovdd.n1340 4.49246
R16305 iovdd.n199 iovdd.n115 4.49246
R16306 iovdd.n1353 iovdd.n1341 4.49246
R16307 iovdd.n202 iovdd.n115 4.49246
R16308 iovdd.n1353 iovdd.n1342 4.49246
R16309 iovdd.n205 iovdd.n115 4.49246
R16310 iovdd.n1353 iovdd.n1343 4.49246
R16311 iovdd.n208 iovdd.n115 4.49246
R16312 iovdd.n1353 iovdd.n1344 4.49246
R16313 iovdd.n211 iovdd.n115 4.49246
R16314 iovdd.n1353 iovdd.n1345 4.49246
R16315 iovdd.n214 iovdd.n115 4.49246
R16316 iovdd.n1353 iovdd.n1346 4.49246
R16317 iovdd.n217 iovdd.n115 4.49246
R16318 iovdd.n1353 iovdd.n1347 4.49246
R16319 iovdd.n220 iovdd.n115 4.49246
R16320 iovdd.n1353 iovdd.n1348 4.49246
R16321 iovdd.n223 iovdd.n115 4.49246
R16322 iovdd.n1353 iovdd.n1349 4.49246
R16323 iovdd.n226 iovdd.n115 4.49246
R16324 iovdd.n1353 iovdd.n1350 4.49246
R16325 iovdd.n229 iovdd.n115 4.49246
R16326 iovdd.n1353 iovdd.n1351 4.49246
R16327 iovdd.n232 iovdd.n115 4.49246
R16328 iovdd.n1353 iovdd.n1352 4.49246
R16329 iovdd.n237 iovdd.n115 4.49246
R16330 iovdd.n1304 iovdd.n401 4.49246
R16331 iovdd.n1298 iovdd.n389 4.49246
R16332 iovdd.n1301 iovdd.n1281 4.49246
R16333 iovdd.n402 iovdd.n389 4.49246
R16334 iovdd.n1301 iovdd.n1280 4.49246
R16335 iovdd.n405 iovdd.n389 4.49246
R16336 iovdd.n1301 iovdd.n1279 4.49246
R16337 iovdd.n408 iovdd.n389 4.49246
R16338 iovdd.n1302 iovdd.n1301 4.49246
R16339 iovdd.n411 iovdd.n389 4.49246
R16340 iovdd.n1301 iovdd.n390 4.49246
R16341 iovdd.n1249 iovdd.n559 4.49246
R16342 iovdd.n1264 iovdd.n560 4.49246
R16343 iovdd.n1252 iovdd.n559 4.49246
R16344 iovdd.n1264 iovdd.n561 4.49246
R16345 iovdd.n1255 iovdd.n559 4.49246
R16346 iovdd.n1264 iovdd.n562 4.49246
R16347 iovdd.n1258 iovdd.n559 4.49246
R16348 iovdd.n1264 iovdd.n563 4.49246
R16349 iovdd.n566 iovdd.n559 4.49246
R16350 iovdd.n1264 iovdd.n1263 4.49246
R16351 iovdd.n564 iovdd.n559 4.49246
R16352 iovdd.n785 iovdd.n774 4.49246
R16353 iovdd.n1236 iovdd.n775 4.49246
R16354 iovdd.n787 iovdd.n774 4.49246
R16355 iovdd.n1236 iovdd.n776 4.49246
R16356 iovdd.n789 iovdd.n774 4.49246
R16357 iovdd.n1236 iovdd.n777 4.49246
R16358 iovdd.n779 iovdd.n774 4.49246
R16359 iovdd.n1236 iovdd.n1235 4.49246
R16360 iovdd.n774 iovdd.n569 4.49246
R16361 iovdd.n1233 iovdd.n568 4.49246
R16362 iovdd.n1236 iovdd.n770 4.49246
R16363 iovdd.n298 iovdd.n272 3.0005
R16364 iovdd.n1262 iovdd.n1240 3.0005
R16365 iovdd.n483 iovdd.n482 3.0005
R16366 iovdd.n474 iovdd.n473 3.0005
R16367 iovdd.n472 iovdd.n471 3.0005
R16368 iovdd.n470 iovdd.n469 3.0005
R16369 iovdd.n468 iovdd.n467 3.0005
R16370 iovdd.n498 iovdd.n497 3.0005
R16371 iovdd.n501 iovdd.n500 3.0005
R16372 iovdd.n504 iovdd.n503 3.0005
R16373 iovdd.n507 iovdd.n506 3.0005
R16374 iovdd.n510 iovdd.n509 3.0005
R16375 iovdd.n458 iovdd.n457 3.0005
R16376 iovdd.n456 iovdd.n455 3.0005
R16377 iovdd.n454 iovdd.n453 3.0005
R16378 iovdd.n452 iovdd.n451 3.0005
R16379 iovdd.n450 iovdd.n449 3.0005
R16380 iovdd.n525 iovdd.n524 3.0005
R16381 iovdd.n528 iovdd.n527 3.0005
R16382 iovdd.n531 iovdd.n530 3.0005
R16383 iovdd.n534 iovdd.n533 3.0005
R16384 iovdd.n440 iovdd.n439 3.0005
R16385 iovdd.n438 iovdd.n437 3.0005
R16386 iovdd.n436 iovdd.n435 3.0005
R16387 iovdd.n434 iovdd.n433 3.0005
R16388 iovdd.n550 iovdd.n549 3.0005
R16389 iovdd.n430 iovdd.n429 3.0005
R16390 iovdd.n556 iovdd.n427 3.0005
R16391 iovdd.n424 iovdd.n423 3.0005
R16392 iovdd.n1248 iovdd.n1247 3.0005
R16393 iovdd.n1254 iovdd.n1253 3.0005
R16394 iovdd.n1257 iovdd.n1256 3.0005
R16395 iovdd.n1260 iovdd.n1259 3.0005
R16396 iovdd.n1242 iovdd.n1241 3.0005
R16397 iovdd.n1244 iovdd.n1243 3.0005
R16398 iovdd.n1246 iovdd.n1245 3.0005
R16399 iovdd.n1251 iovdd.n1250 3.0005
R16400 iovdd.n557 iovdd.n426 3.0005
R16401 iovdd.n555 iovdd.n428 3.0005
R16402 iovdd.n551 iovdd.n432 3.0005
R16403 iovdd.n546 iovdd.n545 3.0005
R16404 iovdd.n543 iovdd.n542 3.0005
R16405 iovdd.n540 iovdd.n539 3.0005
R16406 iovdd.n537 iovdd.n536 3.0005
R16407 iovdd.n442 iovdd.n441 3.0005
R16408 iovdd.n444 iovdd.n443 3.0005
R16409 iovdd.n446 iovdd.n445 3.0005
R16410 iovdd.n448 iovdd.n447 3.0005
R16411 iovdd.n522 iovdd.n521 3.0005
R16412 iovdd.n519 iovdd.n518 3.0005
R16413 iovdd.n516 iovdd.n515 3.0005
R16414 iovdd.n513 iovdd.n512 3.0005
R16415 iovdd.n460 iovdd.n459 3.0005
R16416 iovdd.n462 iovdd.n461 3.0005
R16417 iovdd.n464 iovdd.n463 3.0005
R16418 iovdd.n466 iovdd.n465 3.0005
R16419 iovdd.n495 iovdd.n494 3.0005
R16420 iovdd.n492 iovdd.n491 3.0005
R16421 iovdd.n489 iovdd.n488 3.0005
R16422 iovdd.n486 iovdd.n485 3.0005
R16423 iovdd.n476 iovdd.n475 3.0005
R16424 iovdd.n479 iovdd.n478 3.0005
R16425 iovdd.n300 iovdd.n273 3.0005
R16426 iovdd.n552 iovdd.n551 3.0005
R16427 iovdd.n553 iovdd.n430 3.0005
R16428 iovdd.n555 iovdd.n554 3.0005
R16429 iovdd.n556 iovdd.n425 3.0005
R16430 iovdd.n558 iovdd.n557 3.0005
R16431 iovdd.n1194 iovdd.n1090 3.0005
R16432 iovdd.n1192 iovdd.n1190 3.0005
R16433 iovdd.n1189 iovdd.n1182 3.0005
R16434 iovdd.n1188 iovdd.n1187 3.0005
R16435 iovdd.n1185 iovdd.n1183 3.0005
R16436 iovdd.n1306 iovdd.n387 3.0005
R16437 iovdd.n1306 iovdd.n388 3.0005
R16438 iovdd.n772 iovdd.n565 3.0005
R16439 iovdd.n773 iovdd.n772 3.0005
R16440 iovdd.n862 iovdd.n859 3.0005
R16441 iovdd.n1238 iovdd.n1237 3.0005
R16442 iovdd.n855 iovdd.n778 3.0005
R16443 iovdd.n1234 iovdd.n780 3.0005
R16444 iovdd.n853 iovdd.n782 3.0005
R16445 iovdd.n1232 iovdd.n1231 3.0005
R16446 iovdd.n791 iovdd.n783 3.0005
R16447 iovdd.n851 iovdd.n788 3.0005
R16448 iovdd.n849 iovdd.n784 3.0005
R16449 iovdd.n847 iovdd.n786 3.0005
R16450 iovdd.n845 iovdd.n771 3.0005
R16451 iovdd.n1185 iovdd.n1184 3.0005
R16452 iovdd.n1187 iovdd.n1186 3.0005
R16453 iovdd.n1182 iovdd.n1181 3.0005
R16454 iovdd.n1192 iovdd.n1191 3.0005
R16455 iovdd.n1194 iovdd.n1193 3.0005
R16456 iovdd.n1220 iovdd.n1219 3.0005
R16457 iovdd.n1092 iovdd.n1091 3.0005
R16458 iovdd.n1180 iovdd.n1179 3.0005
R16459 iovdd.n1094 iovdd.n1093 3.0005
R16460 iovdd.n1178 iovdd.n1177 3.0005
R16461 iovdd.n1096 iovdd.n1095 3.0005
R16462 iovdd.n1176 iovdd.n1175 3.0005
R16463 iovdd.n1098 iovdd.n1097 3.0005
R16464 iovdd.n1174 iovdd.n1173 3.0005
R16465 iovdd.n1100 iovdd.n1099 3.0005
R16466 iovdd.n1172 iovdd.n1171 3.0005
R16467 iovdd.n1102 iovdd.n1101 3.0005
R16468 iovdd.n1170 iovdd.n1169 3.0005
R16469 iovdd.n1104 iovdd.n1103 3.0005
R16470 iovdd.n1168 iovdd.n1167 3.0005
R16471 iovdd.n1106 iovdd.n1105 3.0005
R16472 iovdd.n1166 iovdd.n1165 3.0005
R16473 iovdd.n1108 iovdd.n1107 3.0005
R16474 iovdd.n1164 iovdd.n1163 3.0005
R16475 iovdd.n1110 iovdd.n1109 3.0005
R16476 iovdd.n1162 iovdd.n1161 3.0005
R16477 iovdd.n1112 iovdd.n1111 3.0005
R16478 iovdd.n1160 iovdd.n1159 3.0005
R16479 iovdd.n1114 iovdd.n1113 3.0005
R16480 iovdd.n1158 iovdd.n1157 3.0005
R16481 iovdd.n1116 iovdd.n1115 3.0005
R16482 iovdd.n1156 iovdd.n1155 3.0005
R16483 iovdd.n1118 iovdd.n1117 3.0005
R16484 iovdd.n1154 iovdd.n1153 3.0005
R16485 iovdd.n1120 iovdd.n1119 3.0005
R16486 iovdd.n1152 iovdd.n1151 3.0005
R16487 iovdd.n1122 iovdd.n1121 3.0005
R16488 iovdd.n1150 iovdd.n1149 3.0005
R16489 iovdd.n1124 iovdd.n1123 3.0005
R16490 iovdd.n1148 iovdd.n1147 3.0005
R16491 iovdd.n1126 iovdd.n1125 3.0005
R16492 iovdd.n1146 iovdd.n1145 3.0005
R16493 iovdd.n1128 iovdd.n1127 3.0005
R16494 iovdd.n1144 iovdd.n1143 3.0005
R16495 iovdd.n1130 iovdd.n1129 3.0005
R16496 iovdd.n1142 iovdd.n1141 3.0005
R16497 iovdd.n1132 iovdd.n1131 3.0005
R16498 iovdd.n1140 iovdd.n1139 3.0005
R16499 iovdd.n1134 iovdd.n1133 3.0005
R16500 iovdd.n1138 iovdd.n1137 3.0005
R16501 iovdd.n1136 iovdd.n1135 3.0005
R16502 iovdd.n1089 iovdd.n1088 3.0005
R16503 iovdd.n165 iovdd.n112 3.0005
R16504 iovdd.n396 iovdd.n395 3.0005
R16505 iovdd.n407 iovdd.n406 3.0005
R16506 iovdd.n398 iovdd.n397 3.0005
R16507 iovdd.n404 iovdd.n403 3.0005
R16508 iovdd.n400 iovdd.n399 3.0005
R16509 iovdd.n1300 iovdd.n1299 3.0005
R16510 iovdd.n1296 iovdd.n1282 3.0005
R16511 iovdd.n1295 iovdd.n1283 3.0005
R16512 iovdd.n1285 iovdd.n1284 3.0005
R16513 iovdd.n1291 iovdd.n1288 3.0005
R16514 iovdd.n1290 iovdd.n1289 3.0005
R16515 iovdd.n236 iovdd.n235 3.0005
R16516 iovdd.n1354 iovdd.n238 3.0005
R16517 iovdd.n120 iovdd.n119 3.0005
R16518 iovdd.n234 iovdd.n233 3.0005
R16519 iovdd.n122 iovdd.n121 3.0005
R16520 iovdd.n231 iovdd.n230 3.0005
R16521 iovdd.n124 iovdd.n123 3.0005
R16522 iovdd.n228 iovdd.n227 3.0005
R16523 iovdd.n126 iovdd.n125 3.0005
R16524 iovdd.n225 iovdd.n224 3.0005
R16525 iovdd.n128 iovdd.n127 3.0005
R16526 iovdd.n222 iovdd.n221 3.0005
R16527 iovdd.n130 iovdd.n129 3.0005
R16528 iovdd.n219 iovdd.n218 3.0005
R16529 iovdd.n132 iovdd.n131 3.0005
R16530 iovdd.n216 iovdd.n215 3.0005
R16531 iovdd.n134 iovdd.n133 3.0005
R16532 iovdd.n213 iovdd.n212 3.0005
R16533 iovdd.n136 iovdd.n135 3.0005
R16534 iovdd.n210 iovdd.n209 3.0005
R16535 iovdd.n138 iovdd.n137 3.0005
R16536 iovdd.n207 iovdd.n206 3.0005
R16537 iovdd.n140 iovdd.n139 3.0005
R16538 iovdd.n204 iovdd.n203 3.0005
R16539 iovdd.n142 iovdd.n141 3.0005
R16540 iovdd.n201 iovdd.n200 3.0005
R16541 iovdd.n144 iovdd.n143 3.0005
R16542 iovdd.n198 iovdd.n197 3.0005
R16543 iovdd.n146 iovdd.n145 3.0005
R16544 iovdd.n195 iovdd.n194 3.0005
R16545 iovdd.n148 iovdd.n147 3.0005
R16546 iovdd.n192 iovdd.n191 3.0005
R16547 iovdd.n150 iovdd.n149 3.0005
R16548 iovdd.n189 iovdd.n188 3.0005
R16549 iovdd.n152 iovdd.n151 3.0005
R16550 iovdd.n186 iovdd.n185 3.0005
R16551 iovdd.n154 iovdd.n153 3.0005
R16552 iovdd.n183 iovdd.n182 3.0005
R16553 iovdd.n156 iovdd.n155 3.0005
R16554 iovdd.n180 iovdd.n179 3.0005
R16555 iovdd.n158 iovdd.n157 3.0005
R16556 iovdd.n177 iovdd.n176 3.0005
R16557 iovdd.n160 iovdd.n159 3.0005
R16558 iovdd.n174 iovdd.n173 3.0005
R16559 iovdd.n162 iovdd.n161 3.0005
R16560 iovdd.n171 iovdd.n170 3.0005
R16561 iovdd.n164 iovdd.n163 3.0005
R16562 iovdd.n168 iovdd.n167 3.0005
R16563 iovdd.n1303 iovdd.n412 3.0005
R16564 iovdd.n1306 iovdd.n1305 3.0005
R16565 iovdd.n772 iovdd.n392 3.0005
R16566 iovdd.n394 iovdd.n393 3.0005
R16567 iovdd.n410 iovdd.n409 3.0005
R16568 iovdd.n1286 iovdd.n236 3.0005
R16569 iovdd.n1290 iovdd.n1287 3.0005
R16570 iovdd.n1292 iovdd.n1291 3.0005
R16571 iovdd.n1293 iovdd.n1285 3.0005
R16572 iovdd.n1295 iovdd.n1294 3.0005
R16573 iovdd.t0 iovdd.n24 2.83433
R16574 iovdd.t0 iovdd.n21 2.83433
R16575 iovdd.t0 iovdd.n18 2.83433
R16576 iovdd.t0 iovdd.n15 2.83433
R16577 iovdd.t0 iovdd.n2 2.83433
R16578 iovdd.n1361 iovdd.t0 2.83433
R16579 iovdd.t0 iovdd.n6 2.83433
R16580 iovdd.t0 iovdd.n41 2.83433
R16581 iovdd.t0 iovdd.n38 2.83433
R16582 iovdd.t0 iovdd.n35 2.83433
R16583 iovdd.t0 iovdd.n32 2.83433
R16584 iovdd.t0 iovdd.n29 2.83433
R16585 iovdd.t0 iovdd.n26 2.83433
R16586 iovdd.n1309 iovdd.n360 2.82693
R16587 iovdd.n1309 iovdd.n358 2.82693
R16588 iovdd.n1309 iovdd.n355 2.82693
R16589 iovdd.n1309 iovdd.n353 2.82693
R16590 iovdd.n1309 iovdd.n351 2.82693
R16591 iovdd.n1309 iovdd.n349 2.82693
R16592 iovdd.n1309 iovdd.n346 2.82693
R16593 iovdd.n1309 iovdd.n344 2.82693
R16594 iovdd.n1309 iovdd.n342 2.82693
R16595 iovdd.n1309 iovdd.n340 2.82693
R16596 iovdd.n1309 iovdd.n337 2.82693
R16597 iovdd.n1309 iovdd.n335 2.82693
R16598 iovdd.n1309 iovdd.n333 2.82693
R16599 iovdd.n1309 iovdd.n331 2.82693
R16600 iovdd.n1309 iovdd.n328 2.82693
R16601 iovdd.n1309 iovdd.n326 2.82693
R16602 iovdd.n1309 iovdd.n324 2.82693
R16603 iovdd.n1309 iovdd.n321 2.82693
R16604 iovdd.n1309 iovdd.n319 2.82693
R16605 iovdd.n1309 iovdd.n317 2.82693
R16606 iovdd.n1309 iovdd.n315 2.82693
R16607 iovdd.n1309 iovdd.n312 2.82693
R16608 iovdd.n1309 iovdd.n310 2.82693
R16609 iovdd.n1309 iovdd.n308 2.82693
R16610 iovdd.n1309 iovdd.n306 2.82693
R16611 iovdd.n1309 iovdd.n303 2.82693
R16612 iovdd.n1309 iovdd.n301 2.82693
R16613 iovdd.n1229 iovdd.n856 2.82693
R16614 iovdd.n1229 iovdd.n790 2.82693
R16615 iovdd.n1229 iovdd.n850 2.82693
R16616 iovdd.n1229 iovdd.n846 2.82693
R16617 iovdd.n1229 iovdd.n843 2.82693
R16618 iovdd.n1229 iovdd.n841 2.82693
R16619 iovdd.n1229 iovdd.n838 2.82693
R16620 iovdd.n1229 iovdd.n836 2.82693
R16621 iovdd.n1229 iovdd.n834 2.82693
R16622 iovdd.n1229 iovdd.n832 2.82693
R16623 iovdd.n1229 iovdd.n829 2.82693
R16624 iovdd.n1229 iovdd.n827 2.82693
R16625 iovdd.n1229 iovdd.n825 2.82693
R16626 iovdd.n1229 iovdd.n822 2.82693
R16627 iovdd.n1229 iovdd.n820 2.82693
R16628 iovdd.n1229 iovdd.n818 2.82693
R16629 iovdd.n1229 iovdd.n816 2.82693
R16630 iovdd.n1229 iovdd.n813 2.82693
R16631 iovdd.n1229 iovdd.n811 2.82693
R16632 iovdd.n1229 iovdd.n809 2.82693
R16633 iovdd.n1229 iovdd.n807 2.82693
R16634 iovdd.n1229 iovdd.n804 2.82693
R16635 iovdd.n1229 iovdd.n802 2.82693
R16636 iovdd.n1229 iovdd.n800 2.82693
R16637 iovdd.n1229 iovdd.n798 2.82693
R16638 iovdd.n1229 iovdd.n795 2.82693
R16639 iovdd.n1229 iovdd.n793 2.82693
R16640 iovdd.n1359 iovdd.n109 2.82693
R16641 iovdd.n1359 iovdd.n107 2.82693
R16642 iovdd.n1359 iovdd.n104 2.82693
R16643 iovdd.n1359 iovdd.n102 2.82693
R16644 iovdd.n1359 iovdd.n100 2.82693
R16645 iovdd.n1359 iovdd.n98 2.82693
R16646 iovdd.n1359 iovdd.n95 2.82693
R16647 iovdd.n1359 iovdd.n93 2.82693
R16648 iovdd.n1359 iovdd.n91 2.82693
R16649 iovdd.n1359 iovdd.n89 2.82693
R16650 iovdd.n1359 iovdd.n86 2.82693
R16651 iovdd.n1359 iovdd.n84 2.82693
R16652 iovdd.n1359 iovdd.n82 2.82693
R16653 iovdd.n1359 iovdd.n79 2.82693
R16654 iovdd.n1359 iovdd.n77 2.82693
R16655 iovdd.n1359 iovdd.n75 2.82693
R16656 iovdd.n1359 iovdd.n73 2.82693
R16657 iovdd.n1359 iovdd.n70 2.82693
R16658 iovdd.n1359 iovdd.n68 2.82693
R16659 iovdd.n1359 iovdd.n66 2.82693
R16660 iovdd.n1359 iovdd.n64 2.82693
R16661 iovdd.n1359 iovdd.n61 2.82693
R16662 iovdd.n1359 iovdd.n59 2.82693
R16663 iovdd.n1359 iovdd.n57 2.82693
R16664 iovdd.n1359 iovdd.n55 2.82693
R16665 iovdd.n1359 iovdd.n52 2.82693
R16666 iovdd.n1359 iovdd.n50 2.82693
R16667 iovdd.n279 iovdd.n278 2.82693
R16668 iovdd.n281 iovdd.n280 2.82693
R16669 iovdd.n283 iovdd.n282 2.82693
R16670 iovdd.n285 iovdd.n284 2.82693
R16671 iovdd.n287 iovdd.n286 2.82693
R16672 iovdd.n296 iovdd.n291 2.82693
R16673 iovdd.n295 iovdd.n292 2.82693
R16674 iovdd.n294 iovdd.n293 2.82693
R16675 iovdd.n14 iovdd.n1 2.82693
R16676 iovdd.n1363 iovdd.n1362 2.82693
R16677 iovdd.n944 iovdd.n937 0.826084
R16678 iovdd.n649 iovdd.n642 0.826084
R16679 iovdd.n1326 iovdd.n1325 0.822133
R16680 iovdd.n1275 iovdd.n415 0.822133
R16681 iovdd.n943 iovdd.n942 0.818682
R16682 iovdd.n938 iovdd.n936 0.818682
R16683 iovdd.n948 iovdd.n947 0.818682
R16684 iovdd.n949 iovdd.n929 0.818682
R16685 iovdd.n958 iovdd.n957 0.818682
R16686 iovdd.n931 iovdd.n927 0.818682
R16687 iovdd.n963 iovdd.n962 0.818682
R16688 iovdd.n964 iovdd.n920 0.818682
R16689 iovdd.n973 iovdd.n972 0.818682
R16690 iovdd.n922 iovdd.n918 0.818682
R16691 iovdd.n978 iovdd.n977 0.818682
R16692 iovdd.n979 iovdd.n911 0.818682
R16693 iovdd.n988 iovdd.n987 0.818682
R16694 iovdd.n913 iovdd.n909 0.818682
R16695 iovdd.n993 iovdd.n992 0.818682
R16696 iovdd.n994 iovdd.n902 0.818682
R16697 iovdd.n1003 iovdd.n1002 0.818682
R16698 iovdd.n904 iovdd.n900 0.818682
R16699 iovdd.n1008 iovdd.n1007 0.818682
R16700 iovdd.n1009 iovdd.n893 0.818682
R16701 iovdd.n1018 iovdd.n1017 0.818682
R16702 iovdd.n895 iovdd.n891 0.818682
R16703 iovdd.n1023 iovdd.n1022 0.818682
R16704 iovdd.n1024 iovdd.n884 0.818682
R16705 iovdd.n1033 iovdd.n1032 0.818682
R16706 iovdd.n886 iovdd.n882 0.818682
R16707 iovdd.n1038 iovdd.n1037 0.818682
R16708 iovdd.n1039 iovdd.n875 0.818682
R16709 iovdd.n1048 iovdd.n1047 0.818682
R16710 iovdd.n877 iovdd.n873 0.818682
R16711 iovdd.n1053 iovdd.n1052 0.818682
R16712 iovdd.n1054 iovdd.n866 0.818682
R16713 iovdd.n1063 iovdd.n1062 0.818682
R16714 iovdd.n868 iovdd.n246 0.818682
R16715 iovdd.n1316 iovdd.n1315 0.818682
R16716 iovdd.n1318 iovdd.n240 0.818682
R16717 iovdd.n1327 iovdd.n241 0.818682
R16718 iovdd.n1326 iovdd.n118 0.818682
R16719 iovdd.n1328 iovdd.n1327 0.818682
R16720 iovdd.n240 iovdd.n239 0.818682
R16721 iovdd.n1315 iovdd.n1314 0.818682
R16722 iovdd.n247 iovdd.n246 0.818682
R16723 iovdd.n1064 iovdd.n1063 0.818682
R16724 iovdd.n866 iovdd.n865 0.818682
R16725 iovdd.n1052 iovdd.n1051 0.818682
R16726 iovdd.n1050 iovdd.n873 0.818682
R16727 iovdd.n1049 iovdd.n1048 0.818682
R16728 iovdd.n875 iovdd.n874 0.818682
R16729 iovdd.n1037 iovdd.n1036 0.818682
R16730 iovdd.n1035 iovdd.n882 0.818682
R16731 iovdd.n1034 iovdd.n1033 0.818682
R16732 iovdd.n884 iovdd.n883 0.818682
R16733 iovdd.n1022 iovdd.n1021 0.818682
R16734 iovdd.n1020 iovdd.n891 0.818682
R16735 iovdd.n1019 iovdd.n1018 0.818682
R16736 iovdd.n893 iovdd.n892 0.818682
R16737 iovdd.n1007 iovdd.n1006 0.818682
R16738 iovdd.n1005 iovdd.n900 0.818682
R16739 iovdd.n1004 iovdd.n1003 0.818682
R16740 iovdd.n902 iovdd.n901 0.818682
R16741 iovdd.n992 iovdd.n991 0.818682
R16742 iovdd.n990 iovdd.n909 0.818682
R16743 iovdd.n989 iovdd.n988 0.818682
R16744 iovdd.n911 iovdd.n910 0.818682
R16745 iovdd.n977 iovdd.n976 0.818682
R16746 iovdd.n975 iovdd.n918 0.818682
R16747 iovdd.n974 iovdd.n973 0.818682
R16748 iovdd.n920 iovdd.n919 0.818682
R16749 iovdd.n962 iovdd.n961 0.818682
R16750 iovdd.n960 iovdd.n927 0.818682
R16751 iovdd.n959 iovdd.n958 0.818682
R16752 iovdd.n929 iovdd.n928 0.818682
R16753 iovdd.n947 iovdd.n946 0.818682
R16754 iovdd.n945 iovdd.n936 0.818682
R16755 iovdd.n415 iovdd.n391 0.818682
R16756 iovdd.n769 iovdd.n768 0.818682
R16757 iovdd.n571 iovdd.n570 0.818682
R16758 iovdd.n757 iovdd.n756 0.818682
R16759 iovdd.n755 iovdd.n578 0.818682
R16760 iovdd.n754 iovdd.n753 0.818682
R16761 iovdd.n580 iovdd.n579 0.818682
R16762 iovdd.n742 iovdd.n741 0.818682
R16763 iovdd.n740 iovdd.n587 0.818682
R16764 iovdd.n739 iovdd.n738 0.818682
R16765 iovdd.n589 iovdd.n588 0.818682
R16766 iovdd.n727 iovdd.n726 0.818682
R16767 iovdd.n725 iovdd.n596 0.818682
R16768 iovdd.n724 iovdd.n723 0.818682
R16769 iovdd.n598 iovdd.n597 0.818682
R16770 iovdd.n712 iovdd.n711 0.818682
R16771 iovdd.n710 iovdd.n605 0.818682
R16772 iovdd.n709 iovdd.n708 0.818682
R16773 iovdd.n607 iovdd.n606 0.818682
R16774 iovdd.n697 iovdd.n696 0.818682
R16775 iovdd.n695 iovdd.n614 0.818682
R16776 iovdd.n694 iovdd.n693 0.818682
R16777 iovdd.n616 iovdd.n615 0.818682
R16778 iovdd.n682 iovdd.n681 0.818682
R16779 iovdd.n680 iovdd.n623 0.818682
R16780 iovdd.n679 iovdd.n678 0.818682
R16781 iovdd.n625 iovdd.n624 0.818682
R16782 iovdd.n667 iovdd.n666 0.818682
R16783 iovdd.n665 iovdd.n632 0.818682
R16784 iovdd.n664 iovdd.n663 0.818682
R16785 iovdd.n634 iovdd.n633 0.818682
R16786 iovdd.n652 iovdd.n651 0.818682
R16787 iovdd.n650 iovdd.n641 0.818682
R16788 iovdd.n422 iovdd.n421 0.818682
R16789 iovdd.n1266 iovdd.n1265 0.818682
R16790 iovdd.n414 iovdd.n413 0.818682
R16791 iovdd.n1278 iovdd.n1277 0.818682
R16792 iovdd.n648 iovdd.n647 0.818682
R16793 iovdd.n643 iovdd.n641 0.818682
R16794 iovdd.n653 iovdd.n652 0.818682
R16795 iovdd.n654 iovdd.n634 0.818682
R16796 iovdd.n663 iovdd.n662 0.818682
R16797 iovdd.n636 iovdd.n632 0.818682
R16798 iovdd.n668 iovdd.n667 0.818682
R16799 iovdd.n669 iovdd.n625 0.818682
R16800 iovdd.n678 iovdd.n677 0.818682
R16801 iovdd.n627 iovdd.n623 0.818682
R16802 iovdd.n683 iovdd.n682 0.818682
R16803 iovdd.n684 iovdd.n616 0.818682
R16804 iovdd.n693 iovdd.n692 0.818682
R16805 iovdd.n618 iovdd.n614 0.818682
R16806 iovdd.n698 iovdd.n697 0.818682
R16807 iovdd.n699 iovdd.n607 0.818682
R16808 iovdd.n708 iovdd.n707 0.818682
R16809 iovdd.n609 iovdd.n605 0.818682
R16810 iovdd.n713 iovdd.n712 0.818682
R16811 iovdd.n714 iovdd.n598 0.818682
R16812 iovdd.n723 iovdd.n722 0.818682
R16813 iovdd.n600 iovdd.n596 0.818682
R16814 iovdd.n728 iovdd.n727 0.818682
R16815 iovdd.n729 iovdd.n589 0.818682
R16816 iovdd.n738 iovdd.n737 0.818682
R16817 iovdd.n591 iovdd.n587 0.818682
R16818 iovdd.n743 iovdd.n742 0.818682
R16819 iovdd.n744 iovdd.n580 0.818682
R16820 iovdd.n753 iovdd.n752 0.818682
R16821 iovdd.n582 iovdd.n578 0.818682
R16822 iovdd.n758 iovdd.n757 0.818682
R16823 iovdd.n759 iovdd.n571 0.818682
R16824 iovdd.n768 iovdd.n767 0.818682
R16825 iovdd.n573 iovdd.n421 0.818682
R16826 iovdd.n1267 iovdd.n1266 0.818682
R16827 iovdd.n1268 iovdd.n414 0.818682
R16828 iovdd.n1277 iovdd.n1276 0.818682
R16829 iovdd.n945 iovdd.n944 0.416993
R16830 iovdd.n650 iovdd.n649 0.416993
R16831 iovdd.n1239 iovdd 0.341436
R16832 iovdd.n939 iovdd.n937 0.201704
R16833 iovdd.n644 iovdd.n642 0.201704
R16834 iovdd.n1325 iovdd.n1324 0.2005
R16835 iovdd.n1317 iovdd.n242 0.2005
R16836 iovdd.n1320 iovdd.n1319 0.2005
R16837 iovdd.n245 iovdd.n244 0.2005
R16838 iovdd.n1061 iovdd.n1060 0.2005
R16839 iovdd.n869 iovdd.n867 0.2005
R16840 iovdd.n1056 iovdd.n1055 0.2005
R16841 iovdd.n872 iovdd.n871 0.2005
R16842 iovdd.n1046 iovdd.n1045 0.2005
R16843 iovdd.n878 iovdd.n876 0.2005
R16844 iovdd.n1041 iovdd.n1040 0.2005
R16845 iovdd.n881 iovdd.n880 0.2005
R16846 iovdd.n1031 iovdd.n1030 0.2005
R16847 iovdd.n887 iovdd.n885 0.2005
R16848 iovdd.n1026 iovdd.n1025 0.2005
R16849 iovdd.n890 iovdd.n889 0.2005
R16850 iovdd.n1016 iovdd.n1015 0.2005
R16851 iovdd.n896 iovdd.n894 0.2005
R16852 iovdd.n1011 iovdd.n1010 0.2005
R16853 iovdd.n899 iovdd.n898 0.2005
R16854 iovdd.n1001 iovdd.n1000 0.2005
R16855 iovdd.n905 iovdd.n903 0.2005
R16856 iovdd.n996 iovdd.n995 0.2005
R16857 iovdd.n908 iovdd.n907 0.2005
R16858 iovdd.n986 iovdd.n985 0.2005
R16859 iovdd.n914 iovdd.n912 0.2005
R16860 iovdd.n981 iovdd.n980 0.2005
R16861 iovdd.n917 iovdd.n916 0.2005
R16862 iovdd.n971 iovdd.n970 0.2005
R16863 iovdd.n923 iovdd.n921 0.2005
R16864 iovdd.n966 iovdd.n965 0.2005
R16865 iovdd.n926 iovdd.n925 0.2005
R16866 iovdd.n956 iovdd.n955 0.2005
R16867 iovdd.n932 iovdd.n930 0.2005
R16868 iovdd.n951 iovdd.n950 0.2005
R16869 iovdd.n935 iovdd.n934 0.2005
R16870 iovdd.n941 iovdd.n940 0.2005
R16871 iovdd.n1275 iovdd.n1274 0.2005
R16872 iovdd.n417 iovdd.n416 0.2005
R16873 iovdd.n1270 iovdd.n1269 0.2005
R16874 iovdd.n420 iovdd.n419 0.2005
R16875 iovdd.n766 iovdd.n765 0.2005
R16876 iovdd.n574 iovdd.n572 0.2005
R16877 iovdd.n761 iovdd.n760 0.2005
R16878 iovdd.n577 iovdd.n576 0.2005
R16879 iovdd.n751 iovdd.n750 0.2005
R16880 iovdd.n583 iovdd.n581 0.2005
R16881 iovdd.n746 iovdd.n745 0.2005
R16882 iovdd.n586 iovdd.n585 0.2005
R16883 iovdd.n736 iovdd.n735 0.2005
R16884 iovdd.n592 iovdd.n590 0.2005
R16885 iovdd.n731 iovdd.n730 0.2005
R16886 iovdd.n595 iovdd.n594 0.2005
R16887 iovdd.n721 iovdd.n720 0.2005
R16888 iovdd.n601 iovdd.n599 0.2005
R16889 iovdd.n716 iovdd.n715 0.2005
R16890 iovdd.n604 iovdd.n603 0.2005
R16891 iovdd.n706 iovdd.n705 0.2005
R16892 iovdd.n610 iovdd.n608 0.2005
R16893 iovdd.n701 iovdd.n700 0.2005
R16894 iovdd.n613 iovdd.n612 0.2005
R16895 iovdd.n691 iovdd.n690 0.2005
R16896 iovdd.n619 iovdd.n617 0.2005
R16897 iovdd.n686 iovdd.n685 0.2005
R16898 iovdd.n622 iovdd.n621 0.2005
R16899 iovdd.n676 iovdd.n675 0.2005
R16900 iovdd.n628 iovdd.n626 0.2005
R16901 iovdd.n671 iovdd.n670 0.2005
R16902 iovdd.n631 iovdd.n630 0.2005
R16903 iovdd.n661 iovdd.n660 0.2005
R16904 iovdd.n637 iovdd.n635 0.2005
R16905 iovdd.n656 iovdd.n655 0.2005
R16906 iovdd.n640 iovdd.n639 0.2005
R16907 iovdd.n646 iovdd.n645 0.2005
R16908 iovdd.n1357 iovdd 0.1105
R16909 iovdd.n275 iovdd 0.1105
R16910 iovdd.n1227 iovdd 0.1105
R16911 iovdd.n1324 iovdd.n1323 0.1105
R16912 iovdd.n1322 iovdd.n242 0.1105
R16913 iovdd.n1321 iovdd.n1320 0.1105
R16914 iovdd.n244 iovdd.n243 0.1105
R16915 iovdd.n1060 iovdd.n1059 0.1105
R16916 iovdd.n1058 iovdd.n869 0.1105
R16917 iovdd.n1057 iovdd.n1056 0.1105
R16918 iovdd.n871 iovdd.n870 0.1105
R16919 iovdd.n1045 iovdd.n1044 0.1105
R16920 iovdd.n1043 iovdd.n878 0.1105
R16921 iovdd.n1042 iovdd.n1041 0.1105
R16922 iovdd.n880 iovdd.n879 0.1105
R16923 iovdd.n1030 iovdd.n1029 0.1105
R16924 iovdd.n1028 iovdd.n887 0.1105
R16925 iovdd.n1027 iovdd.n1026 0.1105
R16926 iovdd.n889 iovdd.n888 0.1105
R16927 iovdd.n1015 iovdd.n1014 0.1105
R16928 iovdd.n1013 iovdd.n896 0.1105
R16929 iovdd.n1012 iovdd.n1011 0.1105
R16930 iovdd.n898 iovdd.n897 0.1105
R16931 iovdd.n1000 iovdd.n999 0.1105
R16932 iovdd.n998 iovdd.n905 0.1105
R16933 iovdd.n997 iovdd.n996 0.1105
R16934 iovdd.n907 iovdd.n906 0.1105
R16935 iovdd.n985 iovdd.n984 0.1105
R16936 iovdd.n983 iovdd.n914 0.1105
R16937 iovdd.n982 iovdd.n981 0.1105
R16938 iovdd.n916 iovdd.n915 0.1105
R16939 iovdd.n970 iovdd.n969 0.1105
R16940 iovdd.n968 iovdd.n923 0.1105
R16941 iovdd.n967 iovdd.n966 0.1105
R16942 iovdd.n925 iovdd.n924 0.1105
R16943 iovdd.n955 iovdd.n954 0.1105
R16944 iovdd.n953 iovdd.n932 0.1105
R16945 iovdd.n952 iovdd.n951 0.1105
R16946 iovdd.n934 iovdd.n933 0.1105
R16947 iovdd.n1274 iovdd.n1273 0.1105
R16948 iovdd.n1272 iovdd.n417 0.1105
R16949 iovdd.n1271 iovdd.n1270 0.1105
R16950 iovdd.n419 iovdd.n418 0.1105
R16951 iovdd.n765 iovdd.n764 0.1105
R16952 iovdd.n763 iovdd.n574 0.1105
R16953 iovdd.n762 iovdd.n761 0.1105
R16954 iovdd.n576 iovdd.n575 0.1105
R16955 iovdd.n750 iovdd.n749 0.1105
R16956 iovdd.n748 iovdd.n583 0.1105
R16957 iovdd.n747 iovdd.n746 0.1105
R16958 iovdd.n585 iovdd.n584 0.1105
R16959 iovdd.n735 iovdd.n734 0.1105
R16960 iovdd.n733 iovdd.n592 0.1105
R16961 iovdd.n732 iovdd.n731 0.1105
R16962 iovdd.n594 iovdd.n593 0.1105
R16963 iovdd.n720 iovdd.n719 0.1105
R16964 iovdd.n718 iovdd.n601 0.1105
R16965 iovdd.n717 iovdd.n716 0.1105
R16966 iovdd.n603 iovdd.n602 0.1105
R16967 iovdd.n705 iovdd.n704 0.1105
R16968 iovdd.n703 iovdd.n610 0.1105
R16969 iovdd.n702 iovdd.n701 0.1105
R16970 iovdd.n612 iovdd.n611 0.1105
R16971 iovdd.n690 iovdd.n689 0.1105
R16972 iovdd.n688 iovdd.n619 0.1105
R16973 iovdd.n687 iovdd.n686 0.1105
R16974 iovdd.n621 iovdd.n620 0.1105
R16975 iovdd.n675 iovdd.n674 0.1105
R16976 iovdd.n673 iovdd.n628 0.1105
R16977 iovdd.n672 iovdd.n671 0.1105
R16978 iovdd.n630 iovdd.n629 0.1105
R16979 iovdd.n660 iovdd.n659 0.1105
R16980 iovdd.n658 iovdd.n637 0.1105
R16981 iovdd.n657 iovdd.n656 0.1105
R16982 iovdd.n639 iovdd.n638 0.1105
R16983 iovdd.t0 iovdd.n8 0.063271
R16984 iovdd.t0 iovdd.n25 0.0625942
R16985 iovdd.t0 iovdd.n1360 0.0625838
R16986 iovdd.n1363 iovdd.n1 0.0607875
R16987 iovdd.n294 iovdd.n1 0.0607875
R16988 iovdd.n295 iovdd.n294 0.0607875
R16989 iovdd.n296 iovdd.n295 0.0607875
R16990 iovdd.n287 iovdd.n285 0.0607875
R16991 iovdd.n285 iovdd.n283 0.0607875
R16992 iovdd.n283 iovdd.n281 0.0607875
R16993 iovdd.n281 iovdd.n279 0.0607875
R16994 iovdd.n644 iovdd.n638 0.0568704
R16995 iovdd.n939 iovdd.n933 0.0568704
R16996 iovdd iovdd.n1363 0.041993
R16997 iovdd iovdd.n287 0.0350089
R16998 iovdd.n1294 iovdd.n1293 0.0347222
R16999 iovdd.n1293 iovdd.n1292 0.0347222
R17000 iovdd.n1292 iovdd.n1287 0.0347222
R17001 iovdd.n1287 iovdd.n1286 0.0347222
R17002 iovdd.n1188 iovdd.n1183 0.0347222
R17003 iovdd.n1189 iovdd.n1188 0.0347222
R17004 iovdd.n1190 iovdd.n1189 0.0347222
R17005 iovdd.n1190 iovdd.n1090 0.0347222
R17006 iovdd.n558 iovdd.n425 0.0347222
R17007 iovdd.n554 iovdd.n425 0.0347222
R17008 iovdd.n554 iovdd.n553 0.0347222
R17009 iovdd.n553 iovdd.n552 0.0347222
R17010 iovdd.n557 iovdd.n424 0.0347222
R17011 iovdd.n557 iovdd.n556 0.0347222
R17012 iovdd.n556 iovdd.n555 0.0347222
R17013 iovdd.n555 iovdd.n430 0.0347222
R17014 iovdd.n551 iovdd.n430 0.0347222
R17015 iovdd.n551 iovdd.n550 0.0347222
R17016 iovdd.n1185 iovdd.n771 0.0347222
R17017 iovdd.n1187 iovdd.n1185 0.0347222
R17018 iovdd.n1187 iovdd.n1182 0.0347222
R17019 iovdd.n1192 iovdd.n1182 0.0347222
R17020 iovdd.n1194 iovdd.n1192 0.0347222
R17021 iovdd.n1220 iovdd.n1194 0.0347222
R17022 iovdd.n1089 iovdd.n862 0.0347222
R17023 iovdd.n1226 iovdd.n862 0.0347222
R17024 iovdd.n1296 iovdd.n1295 0.0347222
R17025 iovdd.n1295 iovdd.n1285 0.0347222
R17026 iovdd.n1291 iovdd.n1285 0.0347222
R17027 iovdd.n1291 iovdd.n1290 0.0347222
R17028 iovdd.n1290 iovdd.n236 0.0347222
R17029 iovdd.n1354 iovdd.n236 0.0347222
R17030 iovdd.n212 iovdd.n80 0.0301825
R17031 iovdd.n524 iovdd.n330 0.0301825
R17032 iovdd.n1165 iovdd.n823 0.0301825
R17033 iovdd.n1228 iovdd.n858 0.0301825
R17034 iovdd.n45 iovdd.n44 0.0301825
R17035 iovdd.n403 iovdd.n54 0.0293095
R17036 iovdd.n125 iovdd.n71 0.0293095
R17037 iovdd.n143 iovdd.n88 0.0293095
R17038 iovdd.n159 iovdd.n105 0.0293095
R17039 iovdd.n1253 iovdd.n356 0.0293095
R17040 iovdd.n439 iovdd.n339 0.0293095
R17041 iovdd.n457 iovdd.n322 0.0293095
R17042 iovdd.n473 iovdd.n305 0.0293095
R17043 iovdd.n852 iovdd.n851 0.0293095
R17044 iovdd.n1097 iovdd.n831 0.0293095
R17045 iovdd.n1115 iovdd.n814 0.0293095
R17046 iovdd.n1131 iovdd.n797 0.0293095
R17047 iovdd.n133 iovdd.n79 0.0288977
R17048 iovdd.n447 iovdd.n331 0.0288977
R17049 iovdd.n1107 iovdd.n822 0.0288977
R17050 iovdd.n1289 iovdd.n62 0.0284365
R17051 iovdd.n238 iovdd.n63 0.0284365
R17052 iovdd.n188 iovdd.n96 0.0284365
R17053 iovdd.n185 iovdd.n97 0.0284365
R17054 iovdd.n429 iovdd.n348 0.0284365
R17055 iovdd.n549 iovdd.n347 0.0284365
R17056 iovdd.n500 iovdd.n314 0.0284365
R17057 iovdd.n497 iovdd.n313 0.0284365
R17058 iovdd.n1191 iovdd.n840 0.0284365
R17059 iovdd.n1219 iovdd.n839 0.0284365
R17060 iovdd.n1149 iovdd.n806 0.0284365
R17061 iovdd.n1147 iovdd.n805 0.0284365
R17062 iovdd.n1311 iovdd.n1310 0.0284365
R17063 iovdd.n290 iovdd.n277 0.0284365
R17064 iovdd.n399 iovdd.n55 0.0280247
R17065 iovdd.n227 iovdd.n70 0.0280247
R17066 iovdd.n197 iovdd.n89 0.0280247
R17067 iovdd.n176 iovdd.n104 0.0280247
R17068 iovdd.n1247 iovdd.n355 0.0280247
R17069 iovdd.n539 iovdd.n340 0.0280247
R17070 iovdd.n509 iovdd.n321 0.0280247
R17071 iovdd.n488 iovdd.n306 0.0280247
R17072 iovdd.n850 iovdd.n849 0.0280247
R17073 iovdd.n1175 iovdd.n832 0.0280247
R17074 iovdd.n1155 iovdd.n813 0.0280247
R17075 iovdd.n1141 iovdd.n798 0.0280247
R17076 iovdd.n406 iovdd.n53 0.0275635
R17077 iovdd.n127 iovdd.n72 0.0275635
R17078 iovdd.n141 iovdd.n87 0.0275635
R17079 iovdd.n161 iovdd.n106 0.0275635
R17080 iovdd.n1256 iovdd.n357 0.0275635
R17081 iovdd.n441 iovdd.n338 0.0275635
R17082 iovdd.n455 iovdd.n323 0.0275635
R17083 iovdd.n475 iovdd.n304 0.0275635
R17084 iovdd.n1231 iovdd.n1230 0.0275635
R17085 iovdd.n1099 iovdd.n830 0.0275635
R17086 iovdd.n1113 iovdd.n815 0.0275635
R17087 iovdd.n1133 iovdd.n796 0.0275635
R17088 iovdd.n1288 iovdd.n61 0.0271517
R17089 iovdd.n119 iovdd.n64 0.0271517
R17090 iovdd.n149 iovdd.n95 0.0271517
R17091 iovdd.n153 iovdd.n98 0.0271517
R17092 iovdd.n428 iovdd.n349 0.0271517
R17093 iovdd.n433 iovdd.n346 0.0271517
R17094 iovdd.n463 iovdd.n315 0.0271517
R17095 iovdd.n467 iovdd.n312 0.0271517
R17096 iovdd.n1181 iovdd.n841 0.0271517
R17097 iovdd.n1091 iovdd.n838 0.0271517
R17098 iovdd.n1121 iovdd.n807 0.0271517
R17099 iovdd.n1125 iovdd.n804 0.0271517
R17100 iovdd.n215 iovdd.n78 0.0266905
R17101 iovdd.n209 iovdd.n81 0.0266905
R17102 iovdd.n527 iovdd.n332 0.0266905
R17103 iovdd.n521 iovdd.n329 0.0266905
R17104 iovdd.n1167 iovdd.n824 0.0266905
R17105 iovdd.n1163 iovdd.n821 0.0266905
R17106 iovdd.n395 iovdd.n52 0.0262787
R17107 iovdd.n221 iovdd.n73 0.0262787
R17108 iovdd.n203 iovdd.n86 0.0262787
R17109 iovdd.n170 iovdd.n107 0.0262787
R17110 iovdd.n1243 iovdd.n358 0.0262787
R17111 iovdd.n533 iovdd.n337 0.0262787
R17112 iovdd.n515 iovdd.n324 0.0262787
R17113 iovdd.n482 iovdd.n303 0.0262787
R17114 iovdd.n853 iovdd.n790 0.0262787
R17115 iovdd.n1171 iovdd.n829 0.0262787
R17116 iovdd.n1159 iovdd.n816 0.0262787
R17117 iovdd.n1137 iovdd.n795 0.0262787
R17118 iovdd.n1299 iovdd.n56 0.0258175
R17119 iovdd.n123 iovdd.n69 0.0258175
R17120 iovdd.n145 iovdd.n90 0.0258175
R17121 iovdd.n157 iovdd.n103 0.0258175
R17122 iovdd.n1250 iovdd.n354 0.0258175
R17123 iovdd.n437 iovdd.n341 0.0258175
R17124 iovdd.n459 iovdd.n320 0.0258175
R17125 iovdd.n471 iovdd.n307 0.0258175
R17126 iovdd.n848 iovdd.n847 0.0258175
R17127 iovdd.n1095 iovdd.n833 0.0258175
R17128 iovdd.n1117 iovdd.n812 0.0258175
R17129 iovdd.n1129 iovdd.n799 0.0258175
R17130 iovdd.n131 iovdd.n77 0.0254057
R17131 iovdd.n137 iovdd.n82 0.0254057
R17132 iovdd.n445 iovdd.n333 0.0254057
R17133 iovdd.n451 iovdd.n328 0.0254057
R17134 iovdd.n1103 iovdd.n825 0.0254057
R17135 iovdd.n1109 iovdd.n820 0.0254057
R17136 iovdd.n1284 iovdd.n60 0.0249444
R17137 iovdd.n233 iovdd.n65 0.0249444
R17138 iovdd.n191 iovdd.n94 0.0249444
R17139 iovdd.n182 iovdd.n99 0.0249444
R17140 iovdd.n427 iovdd.n350 0.0249444
R17141 iovdd.n545 iovdd.n345 0.0249444
R17142 iovdd.n503 iovdd.n316 0.0249444
R17143 iovdd.n494 iovdd.n311 0.0249444
R17144 iovdd.n1186 iovdd.n842 0.0249444
R17145 iovdd.n1179 iovdd.n837 0.0249444
R17146 iovdd.n1151 iovdd.n808 0.0249444
R17147 iovdd.n1145 iovdd.n803 0.0249444
R17148 iovdd.n1282 iovdd.n57 0.0245327
R17149 iovdd.n230 iovdd.n68 0.0245327
R17150 iovdd.n194 iovdd.n91 0.0245327
R17151 iovdd.n179 iovdd.n102 0.0245327
R17152 iovdd.n423 iovdd.n353 0.0245327
R17153 iovdd.n542 iovdd.n342 0.0245327
R17154 iovdd.n506 iovdd.n319 0.0245327
R17155 iovdd.n491 iovdd.n308 0.0245327
R17156 iovdd.n846 iovdd.n845 0.0245327
R17157 iovdd.n1177 iovdd.n834 0.0245327
R17158 iovdd.n1153 iovdd.n811 0.0245327
R17159 iovdd.n1143 iovdd.n800 0.0245327
R17160 iovdd.n279 iovdd.n111 0.0245327
R17161 iovdd.n409 iovdd.n51 0.0240714
R17162 iovdd.n129 iovdd.n74 0.0240714
R17163 iovdd.n139 iovdd.n85 0.0240714
R17164 iovdd.n163 iovdd.n108 0.0240714
R17165 iovdd.n1259 iovdd.n359 0.0240714
R17166 iovdd.n443 iovdd.n336 0.0240714
R17167 iovdd.n453 iovdd.n325 0.0240714
R17168 iovdd.n478 iovdd.n302 0.0240714
R17169 iovdd.n854 iovdd.n780 0.0240714
R17170 iovdd.n1101 iovdd.n828 0.0240714
R17171 iovdd.n1111 iovdd.n817 0.0240714
R17172 iovdd.n1135 iovdd.n794 0.0240714
R17173 iovdd.n1283 iovdd.n59 0.0236596
R17174 iovdd.n121 iovdd.n66 0.0236596
R17175 iovdd.n147 iovdd.n93 0.0236596
R17176 iovdd.n155 iovdd.n100 0.0236596
R17177 iovdd.n426 iovdd.n351 0.0236596
R17178 iovdd.n435 iovdd.n344 0.0236596
R17179 iovdd.n461 iovdd.n317 0.0236596
R17180 iovdd.n469 iovdd.n310 0.0236596
R17181 iovdd.n1184 iovdd.n843 0.0236596
R17182 iovdd.n1093 iovdd.n836 0.0236596
R17183 iovdd.n1119 iovdd.n809 0.0236596
R17184 iovdd.n1127 iovdd.n802 0.0236596
R17185 iovdd.n393 iovdd.n46 0.0231984
R17186 iovdd.n218 iovdd.n76 0.0231984
R17187 iovdd.n206 iovdd.n83 0.0231984
R17188 iovdd.n167 iovdd.n110 0.0231984
R17189 iovdd.n1241 iovdd.n361 0.0231984
R17190 iovdd.n530 iovdd.n334 0.0231984
R17191 iovdd.n518 iovdd.n327 0.0231984
R17192 iovdd.n300 iovdd.n299 0.0231984
R17193 iovdd.n855 iovdd.n567 0.0231984
R17194 iovdd.n1169 iovdd.n826 0.0231984
R17195 iovdd.n1161 iovdd.n819 0.0231984
R17196 iovdd.n1088 iovdd.n792 0.0231984
R17197 iovdd.n393 iovdd.n50 0.0227866
R17198 iovdd.n218 iovdd.n75 0.0227866
R17199 iovdd.n206 iovdd.n84 0.0227866
R17200 iovdd.n167 iovdd.n109 0.0227866
R17201 iovdd.n1241 iovdd.n360 0.0227866
R17202 iovdd.n530 iovdd.n335 0.0227866
R17203 iovdd.n518 iovdd.n326 0.0227866
R17204 iovdd.n301 iovdd.n300 0.0227866
R17205 iovdd.n856 iovdd.n855 0.0227866
R17206 iovdd.n1169 iovdd.n827 0.0227866
R17207 iovdd.n1161 iovdd.n818 0.0227866
R17208 iovdd.n1088 iovdd.n793 0.0227866
R17209 iovdd.n1283 iovdd.n58 0.0223254
R17210 iovdd.n121 iovdd.n67 0.0223254
R17211 iovdd.n147 iovdd.n92 0.0223254
R17212 iovdd.n155 iovdd.n101 0.0223254
R17213 iovdd.n426 iovdd.n352 0.0223254
R17214 iovdd.n435 iovdd.n343 0.0223254
R17215 iovdd.n461 iovdd.n318 0.0223254
R17216 iovdd.n469 iovdd.n309 0.0223254
R17217 iovdd.n1184 iovdd.n844 0.0223254
R17218 iovdd.n1093 iovdd.n835 0.0223254
R17219 iovdd.n1119 iovdd.n810 0.0223254
R17220 iovdd.n1127 iovdd.n801 0.0223254
R17221 iovdd.n1227 iovdd.n861 0.0223254
R17222 iovdd.n1358 iovdd.n1357 0.0223254
R17223 iovdd.n409 iovdd.n50 0.0219136
R17224 iovdd.n129 iovdd.n75 0.0219136
R17225 iovdd.n139 iovdd.n84 0.0219136
R17226 iovdd.n163 iovdd.n109 0.0219136
R17227 iovdd.n1259 iovdd.n360 0.0219136
R17228 iovdd.n443 iovdd.n335 0.0219136
R17229 iovdd.n453 iovdd.n326 0.0219136
R17230 iovdd.n478 iovdd.n301 0.0219136
R17231 iovdd.n856 iovdd.n780 0.0219136
R17232 iovdd.n1101 iovdd.n827 0.0219136
R17233 iovdd.n1111 iovdd.n818 0.0219136
R17234 iovdd.n1135 iovdd.n793 0.0219136
R17235 iovdd.n1282 iovdd.n58 0.0214524
R17236 iovdd.n230 iovdd.n67 0.0214524
R17237 iovdd.n194 iovdd.n92 0.0214524
R17238 iovdd.n179 iovdd.n101 0.0214524
R17239 iovdd.n423 iovdd.n352 0.0214524
R17240 iovdd.n542 iovdd.n343 0.0214524
R17241 iovdd.n506 iovdd.n318 0.0214524
R17242 iovdd.n491 iovdd.n309 0.0214524
R17243 iovdd.n845 iovdd.n844 0.0214524
R17244 iovdd.n1177 iovdd.n835 0.0214524
R17245 iovdd.n1153 iovdd.n810 0.0214524
R17246 iovdd.n1143 iovdd.n801 0.0214524
R17247 iovdd.n1225 iovdd.n861 0.0214524
R17248 iovdd.n1358 iovdd.n111 0.0214524
R17249 iovdd.n1284 iovdd.n59 0.0210406
R17250 iovdd.n233 iovdd.n66 0.0210406
R17251 iovdd.n191 iovdd.n93 0.0210406
R17252 iovdd.n182 iovdd.n100 0.0210406
R17253 iovdd.n427 iovdd.n351 0.0210406
R17254 iovdd.n545 iovdd.n344 0.0210406
R17255 iovdd.n503 iovdd.n317 0.0210406
R17256 iovdd.n494 iovdd.n310 0.0210406
R17257 iovdd.n1186 iovdd.n843 0.0210406
R17258 iovdd.n1179 iovdd.n836 0.0210406
R17259 iovdd.n1151 iovdd.n809 0.0210406
R17260 iovdd.n1145 iovdd.n802 0.0210406
R17261 iovdd.n412 iovdd.n46 0.0205794
R17262 iovdd.n131 iovdd.n76 0.0205794
R17263 iovdd.n137 iovdd.n83 0.0205794
R17264 iovdd.n112 iovdd.n110 0.0205794
R17265 iovdd.n1240 iovdd.n361 0.0205794
R17266 iovdd.n445 iovdd.n334 0.0205794
R17267 iovdd.n451 iovdd.n327 0.0205794
R17268 iovdd.n299 iovdd.n298 0.0205794
R17269 iovdd.n1238 iovdd.n567 0.0205794
R17270 iovdd.n1103 iovdd.n826 0.0205794
R17271 iovdd.n1109 iovdd.n819 0.0205794
R17272 iovdd.n859 iovdd.n792 0.0205794
R17273 iovdd.n1299 iovdd.n57 0.0201676
R17274 iovdd.n123 iovdd.n68 0.0201676
R17275 iovdd.n145 iovdd.n91 0.0201676
R17276 iovdd.n157 iovdd.n102 0.0201676
R17277 iovdd.n1250 iovdd.n353 0.0201676
R17278 iovdd.n437 iovdd.n342 0.0201676
R17279 iovdd.n459 iovdd.n319 0.0201676
R17280 iovdd.n471 iovdd.n308 0.0201676
R17281 iovdd.n847 iovdd.n846 0.0201676
R17282 iovdd.n1095 iovdd.n834 0.0201676
R17283 iovdd.n1117 iovdd.n811 0.0201676
R17284 iovdd.n1129 iovdd.n800 0.0201676
R17285 iovdd.n395 iovdd.n51 0.0197063
R17286 iovdd.n221 iovdd.n74 0.0197063
R17287 iovdd.n203 iovdd.n85 0.0197063
R17288 iovdd.n170 iovdd.n108 0.0197063
R17289 iovdd.n1243 iovdd.n359 0.0197063
R17290 iovdd.n533 iovdd.n336 0.0197063
R17291 iovdd.n515 iovdd.n325 0.0197063
R17292 iovdd.n482 iovdd.n302 0.0197063
R17293 iovdd.n854 iovdd.n853 0.0197063
R17294 iovdd.n1171 iovdd.n828 0.0197063
R17295 iovdd.n1159 iovdd.n817 0.0197063
R17296 iovdd.n1137 iovdd.n794 0.0197063
R17297 iovdd.n215 iovdd.n77 0.0192946
R17298 iovdd.n209 iovdd.n82 0.0192946
R17299 iovdd.n527 iovdd.n333 0.0192946
R17300 iovdd.n521 iovdd.n328 0.0192946
R17301 iovdd.n1167 iovdd.n825 0.0192946
R17302 iovdd.n1163 iovdd.n820 0.0192946
R17303 iovdd.n1288 iovdd.n60 0.0188333
R17304 iovdd.n119 iovdd.n65 0.0188333
R17305 iovdd.n149 iovdd.n94 0.0188333
R17306 iovdd.n153 iovdd.n99 0.0188333
R17307 iovdd.n428 iovdd.n350 0.0188333
R17308 iovdd.n433 iovdd.n345 0.0188333
R17309 iovdd.n463 iovdd.n316 0.0188333
R17310 iovdd.n467 iovdd.n311 0.0188333
R17311 iovdd.n1181 iovdd.n842 0.0188333
R17312 iovdd.n1091 iovdd.n837 0.0188333
R17313 iovdd.n1121 iovdd.n808 0.0188333
R17314 iovdd.n1125 iovdd.n803 0.0188333
R17315 iovdd.n406 iovdd.n52 0.0184215
R17316 iovdd.n127 iovdd.n73 0.0184215
R17317 iovdd.n141 iovdd.n86 0.0184215
R17318 iovdd.n161 iovdd.n107 0.0184215
R17319 iovdd.n1256 iovdd.n358 0.0184215
R17320 iovdd.n441 iovdd.n337 0.0184215
R17321 iovdd.n455 iovdd.n324 0.0184215
R17322 iovdd.n475 iovdd.n303 0.0184215
R17323 iovdd.n1231 iovdd.n790 0.0184215
R17324 iovdd.n1099 iovdd.n829 0.0184215
R17325 iovdd.n1113 iovdd.n816 0.0184215
R17326 iovdd.n1133 iovdd.n795 0.0184215
R17327 iovdd.n565 iovdd.n564 0.0180786
R17328 iovdd.n1263 iovdd.n1262 0.0180786
R17329 iovdd.n1242 iovdd.n566 0.0180786
R17330 iovdd.n1260 iovdd.n563 0.0180786
R17331 iovdd.n1258 iovdd.n1244 0.0180786
R17332 iovdd.n1257 iovdd.n562 0.0180786
R17333 iovdd.n1255 iovdd.n1246 0.0180786
R17334 iovdd.n1254 iovdd.n561 0.0180786
R17335 iovdd.n1252 iovdd.n1248 0.0180786
R17336 iovdd.n1251 iovdd.n560 0.0180786
R17337 iovdd.n1249 iovdd.n424 0.0180786
R17338 iovdd.n434 iovdd.n249 0.0180786
R17339 iovdd.n546 iovdd.n544 0.0180786
R17340 iovdd.n436 iovdd.n250 0.0180786
R17341 iovdd.n543 iovdd.n541 0.0180786
R17342 iovdd.n438 iovdd.n251 0.0180786
R17343 iovdd.n540 iovdd.n538 0.0180786
R17344 iovdd.n440 iovdd.n252 0.0180786
R17345 iovdd.n537 iovdd.n535 0.0180786
R17346 iovdd.n442 iovdd.n253 0.0180786
R17347 iovdd.n534 iovdd.n532 0.0180786
R17348 iovdd.n444 iovdd.n254 0.0180786
R17349 iovdd.n531 iovdd.n529 0.0180786
R17350 iovdd.n446 iovdd.n255 0.0180786
R17351 iovdd.n528 iovdd.n526 0.0180786
R17352 iovdd.n448 iovdd.n256 0.0180786
R17353 iovdd.n525 iovdd.n523 0.0180786
R17354 iovdd.n450 iovdd.n257 0.0180786
R17355 iovdd.n522 iovdd.n520 0.0180786
R17356 iovdd.n452 iovdd.n258 0.0180786
R17357 iovdd.n519 iovdd.n517 0.0180786
R17358 iovdd.n454 iovdd.n259 0.0180786
R17359 iovdd.n516 iovdd.n514 0.0180786
R17360 iovdd.n456 iovdd.n260 0.0180786
R17361 iovdd.n513 iovdd.n511 0.0180786
R17362 iovdd.n458 iovdd.n261 0.0180786
R17363 iovdd.n510 iovdd.n508 0.0180786
R17364 iovdd.n460 iovdd.n262 0.0180786
R17365 iovdd.n507 iovdd.n505 0.0180786
R17366 iovdd.n462 iovdd.n263 0.0180786
R17367 iovdd.n504 iovdd.n502 0.0180786
R17368 iovdd.n464 iovdd.n264 0.0180786
R17369 iovdd.n501 iovdd.n499 0.0180786
R17370 iovdd.n466 iovdd.n265 0.0180786
R17371 iovdd.n498 iovdd.n496 0.0180786
R17372 iovdd.n468 iovdd.n266 0.0180786
R17373 iovdd.n495 iovdd.n493 0.0180786
R17374 iovdd.n470 iovdd.n267 0.0180786
R17375 iovdd.n492 iovdd.n490 0.0180786
R17376 iovdd.n472 iovdd.n268 0.0180786
R17377 iovdd.n489 iovdd.n487 0.0180786
R17378 iovdd.n474 iovdd.n269 0.0180786
R17379 iovdd.n486 iovdd.n484 0.0180786
R17380 iovdd.n476 iovdd.n270 0.0180786
R17381 iovdd.n483 iovdd.n481 0.0180786
R17382 iovdd.n479 iovdd.n271 0.0180786
R17383 iovdd.n477 iovdd.n273 0.0180786
R17384 iovdd.n480 iovdd.n272 0.0180786
R17385 iovdd.n1312 iovdd.n274 0.0180786
R17386 iovdd.n1312 iovdd.n276 0.0180786
R17387 iovdd.n274 iovdd.n272 0.0180786
R17388 iovdd.n480 iovdd.n273 0.0180786
R17389 iovdd.n479 iovdd.n477 0.0180786
R17390 iovdd.n483 iovdd.n271 0.0180786
R17391 iovdd.n481 iovdd.n476 0.0180786
R17392 iovdd.n486 iovdd.n270 0.0180786
R17393 iovdd.n484 iovdd.n474 0.0180786
R17394 iovdd.n489 iovdd.n269 0.0180786
R17395 iovdd.n487 iovdd.n472 0.0180786
R17396 iovdd.n492 iovdd.n268 0.0180786
R17397 iovdd.n490 iovdd.n470 0.0180786
R17398 iovdd.n495 iovdd.n267 0.0180786
R17399 iovdd.n493 iovdd.n468 0.0180786
R17400 iovdd.n498 iovdd.n266 0.0180786
R17401 iovdd.n496 iovdd.n466 0.0180786
R17402 iovdd.n501 iovdd.n265 0.0180786
R17403 iovdd.n499 iovdd.n464 0.0180786
R17404 iovdd.n504 iovdd.n264 0.0180786
R17405 iovdd.n502 iovdd.n462 0.0180786
R17406 iovdd.n507 iovdd.n263 0.0180786
R17407 iovdd.n505 iovdd.n460 0.0180786
R17408 iovdd.n510 iovdd.n262 0.0180786
R17409 iovdd.n508 iovdd.n458 0.0180786
R17410 iovdd.n513 iovdd.n261 0.0180786
R17411 iovdd.n511 iovdd.n456 0.0180786
R17412 iovdd.n516 iovdd.n260 0.0180786
R17413 iovdd.n514 iovdd.n454 0.0180786
R17414 iovdd.n519 iovdd.n259 0.0180786
R17415 iovdd.n517 iovdd.n452 0.0180786
R17416 iovdd.n522 iovdd.n258 0.0180786
R17417 iovdd.n520 iovdd.n450 0.0180786
R17418 iovdd.n525 iovdd.n257 0.0180786
R17419 iovdd.n523 iovdd.n448 0.0180786
R17420 iovdd.n528 iovdd.n256 0.0180786
R17421 iovdd.n526 iovdd.n446 0.0180786
R17422 iovdd.n531 iovdd.n255 0.0180786
R17423 iovdd.n529 iovdd.n444 0.0180786
R17424 iovdd.n534 iovdd.n254 0.0180786
R17425 iovdd.n532 iovdd.n442 0.0180786
R17426 iovdd.n537 iovdd.n253 0.0180786
R17427 iovdd.n535 iovdd.n440 0.0180786
R17428 iovdd.n540 iovdd.n252 0.0180786
R17429 iovdd.n538 iovdd.n438 0.0180786
R17430 iovdd.n543 iovdd.n251 0.0180786
R17431 iovdd.n541 iovdd.n436 0.0180786
R17432 iovdd.n546 iovdd.n250 0.0180786
R17433 iovdd.n544 iovdd.n434 0.0180786
R17434 iovdd.n550 iovdd.n249 0.0180786
R17435 iovdd.n297 iovdd.n276 0.0180786
R17436 iovdd.n773 iovdd.n770 0.0180786
R17437 iovdd.n1237 iovdd.n568 0.0180786
R17438 iovdd.n778 iovdd.n569 0.0180786
R17439 iovdd.n1235 iovdd.n1234 0.0180786
R17440 iovdd.n782 iovdd.n779 0.0180786
R17441 iovdd.n1232 iovdd.n777 0.0180786
R17442 iovdd.n789 iovdd.n783 0.0180786
R17443 iovdd.n788 iovdd.n776 0.0180786
R17444 iovdd.n787 iovdd.n784 0.0180786
R17445 iovdd.n786 iovdd.n775 0.0180786
R17446 iovdd.n785 iovdd.n771 0.0180786
R17447 iovdd.n1220 iovdd.n1065 0.0180786
R17448 iovdd.n1195 iovdd.n1092 0.0180786
R17449 iovdd.n1180 iovdd.n1066 0.0180786
R17450 iovdd.n1196 iovdd.n1094 0.0180786
R17451 iovdd.n1178 iovdd.n1067 0.0180786
R17452 iovdd.n1197 iovdd.n1096 0.0180786
R17453 iovdd.n1176 iovdd.n1068 0.0180786
R17454 iovdd.n1198 iovdd.n1098 0.0180786
R17455 iovdd.n1174 iovdd.n1069 0.0180786
R17456 iovdd.n1199 iovdd.n1100 0.0180786
R17457 iovdd.n1172 iovdd.n1070 0.0180786
R17458 iovdd.n1200 iovdd.n1102 0.0180786
R17459 iovdd.n1170 iovdd.n1071 0.0180786
R17460 iovdd.n1201 iovdd.n1104 0.0180786
R17461 iovdd.n1168 iovdd.n1072 0.0180786
R17462 iovdd.n1202 iovdd.n1106 0.0180786
R17463 iovdd.n1166 iovdd.n1073 0.0180786
R17464 iovdd.n1203 iovdd.n1108 0.0180786
R17465 iovdd.n1164 iovdd.n1074 0.0180786
R17466 iovdd.n1204 iovdd.n1110 0.0180786
R17467 iovdd.n1162 iovdd.n1075 0.0180786
R17468 iovdd.n1205 iovdd.n1112 0.0180786
R17469 iovdd.n1160 iovdd.n1076 0.0180786
R17470 iovdd.n1206 iovdd.n1114 0.0180786
R17471 iovdd.n1158 iovdd.n1077 0.0180786
R17472 iovdd.n1207 iovdd.n1116 0.0180786
R17473 iovdd.n1156 iovdd.n1078 0.0180786
R17474 iovdd.n1208 iovdd.n1118 0.0180786
R17475 iovdd.n1154 iovdd.n1079 0.0180786
R17476 iovdd.n1209 iovdd.n1120 0.0180786
R17477 iovdd.n1152 iovdd.n1080 0.0180786
R17478 iovdd.n1210 iovdd.n1122 0.0180786
R17479 iovdd.n1150 iovdd.n1081 0.0180786
R17480 iovdd.n1211 iovdd.n1124 0.0180786
R17481 iovdd.n1148 iovdd.n1082 0.0180786
R17482 iovdd.n1212 iovdd.n1126 0.0180786
R17483 iovdd.n1146 iovdd.n1083 0.0180786
R17484 iovdd.n1213 iovdd.n1128 0.0180786
R17485 iovdd.n1144 iovdd.n1084 0.0180786
R17486 iovdd.n1214 iovdd.n1130 0.0180786
R17487 iovdd.n1142 iovdd.n1085 0.0180786
R17488 iovdd.n1215 iovdd.n1132 0.0180786
R17489 iovdd.n1140 iovdd.n1086 0.0180786
R17490 iovdd.n1216 iovdd.n1134 0.0180786
R17491 iovdd.n1138 iovdd.n1087 0.0180786
R17492 iovdd.n1217 iovdd.n1136 0.0180786
R17493 iovdd.n1226 iovdd.n1224 0.0180786
R17494 iovdd.n1217 iovdd.n1089 0.0180786
R17495 iovdd.n1136 iovdd.n1087 0.0180786
R17496 iovdd.n1216 iovdd.n1138 0.0180786
R17497 iovdd.n1134 iovdd.n1086 0.0180786
R17498 iovdd.n1215 iovdd.n1140 0.0180786
R17499 iovdd.n1132 iovdd.n1085 0.0180786
R17500 iovdd.n1214 iovdd.n1142 0.0180786
R17501 iovdd.n1130 iovdd.n1084 0.0180786
R17502 iovdd.n1213 iovdd.n1144 0.0180786
R17503 iovdd.n1128 iovdd.n1083 0.0180786
R17504 iovdd.n1212 iovdd.n1146 0.0180786
R17505 iovdd.n1126 iovdd.n1082 0.0180786
R17506 iovdd.n1211 iovdd.n1148 0.0180786
R17507 iovdd.n1124 iovdd.n1081 0.0180786
R17508 iovdd.n1210 iovdd.n1150 0.0180786
R17509 iovdd.n1122 iovdd.n1080 0.0180786
R17510 iovdd.n1209 iovdd.n1152 0.0180786
R17511 iovdd.n1120 iovdd.n1079 0.0180786
R17512 iovdd.n1208 iovdd.n1154 0.0180786
R17513 iovdd.n1118 iovdd.n1078 0.0180786
R17514 iovdd.n1207 iovdd.n1156 0.0180786
R17515 iovdd.n1116 iovdd.n1077 0.0180786
R17516 iovdd.n1206 iovdd.n1158 0.0180786
R17517 iovdd.n1114 iovdd.n1076 0.0180786
R17518 iovdd.n1205 iovdd.n1160 0.0180786
R17519 iovdd.n1112 iovdd.n1075 0.0180786
R17520 iovdd.n1204 iovdd.n1162 0.0180786
R17521 iovdd.n1110 iovdd.n1074 0.0180786
R17522 iovdd.n1203 iovdd.n1164 0.0180786
R17523 iovdd.n1108 iovdd.n1073 0.0180786
R17524 iovdd.n1202 iovdd.n1166 0.0180786
R17525 iovdd.n1106 iovdd.n1072 0.0180786
R17526 iovdd.n1201 iovdd.n1168 0.0180786
R17527 iovdd.n1104 iovdd.n1071 0.0180786
R17528 iovdd.n1200 iovdd.n1170 0.0180786
R17529 iovdd.n1102 iovdd.n1070 0.0180786
R17530 iovdd.n1199 iovdd.n1172 0.0180786
R17531 iovdd.n1100 iovdd.n1069 0.0180786
R17532 iovdd.n1198 iovdd.n1174 0.0180786
R17533 iovdd.n1098 iovdd.n1068 0.0180786
R17534 iovdd.n1197 iovdd.n1176 0.0180786
R17535 iovdd.n1096 iovdd.n1067 0.0180786
R17536 iovdd.n1196 iovdd.n1178 0.0180786
R17537 iovdd.n1094 iovdd.n1066 0.0180786
R17538 iovdd.n1195 iovdd.n1180 0.0180786
R17539 iovdd.n1092 iovdd.n1065 0.0180786
R17540 iovdd.n1224 iovdd.n860 0.0180786
R17541 iovdd.n392 iovdd.n390 0.0180786
R17542 iovdd.n1303 iovdd.n411 0.0180786
R17543 iovdd.n1302 iovdd.n394 0.0180786
R17544 iovdd.n410 iovdd.n408 0.0180786
R17545 iovdd.n1279 iovdd.n396 0.0180786
R17546 iovdd.n407 iovdd.n405 0.0180786
R17547 iovdd.n1280 iovdd.n398 0.0180786
R17548 iovdd.n404 iovdd.n402 0.0180786
R17549 iovdd.n1281 iovdd.n400 0.0180786
R17550 iovdd.n1300 iovdd.n1298 0.0180786
R17551 iovdd.n1296 iovdd.n401 0.0180786
R17552 iovdd.n237 iovdd.n120 0.0180786
R17553 iovdd.n1352 iovdd.n234 0.0180786
R17554 iovdd.n232 iovdd.n122 0.0180786
R17555 iovdd.n1351 iovdd.n231 0.0180786
R17556 iovdd.n229 iovdd.n124 0.0180786
R17557 iovdd.n1350 iovdd.n228 0.0180786
R17558 iovdd.n226 iovdd.n126 0.0180786
R17559 iovdd.n1349 iovdd.n225 0.0180786
R17560 iovdd.n223 iovdd.n128 0.0180786
R17561 iovdd.n1348 iovdd.n222 0.0180786
R17562 iovdd.n220 iovdd.n130 0.0180786
R17563 iovdd.n1347 iovdd.n219 0.0180786
R17564 iovdd.n217 iovdd.n132 0.0180786
R17565 iovdd.n1346 iovdd.n216 0.0180786
R17566 iovdd.n214 iovdd.n134 0.0180786
R17567 iovdd.n1345 iovdd.n213 0.0180786
R17568 iovdd.n211 iovdd.n136 0.0180786
R17569 iovdd.n1344 iovdd.n210 0.0180786
R17570 iovdd.n208 iovdd.n138 0.0180786
R17571 iovdd.n1343 iovdd.n207 0.0180786
R17572 iovdd.n205 iovdd.n140 0.0180786
R17573 iovdd.n1342 iovdd.n204 0.0180786
R17574 iovdd.n202 iovdd.n142 0.0180786
R17575 iovdd.n1341 iovdd.n201 0.0180786
R17576 iovdd.n199 iovdd.n144 0.0180786
R17577 iovdd.n1340 iovdd.n198 0.0180786
R17578 iovdd.n196 iovdd.n146 0.0180786
R17579 iovdd.n1339 iovdd.n195 0.0180786
R17580 iovdd.n193 iovdd.n148 0.0180786
R17581 iovdd.n1338 iovdd.n192 0.0180786
R17582 iovdd.n190 iovdd.n150 0.0180786
R17583 iovdd.n1337 iovdd.n189 0.0180786
R17584 iovdd.n187 iovdd.n152 0.0180786
R17585 iovdd.n1336 iovdd.n186 0.0180786
R17586 iovdd.n184 iovdd.n154 0.0180786
R17587 iovdd.n1335 iovdd.n183 0.0180786
R17588 iovdd.n181 iovdd.n156 0.0180786
R17589 iovdd.n1334 iovdd.n180 0.0180786
R17590 iovdd.n178 iovdd.n158 0.0180786
R17591 iovdd.n1333 iovdd.n177 0.0180786
R17592 iovdd.n175 iovdd.n160 0.0180786
R17593 iovdd.n1332 iovdd.n174 0.0180786
R17594 iovdd.n172 iovdd.n162 0.0180786
R17595 iovdd.n1331 iovdd.n171 0.0180786
R17596 iovdd.n169 iovdd.n164 0.0180786
R17597 iovdd.n1330 iovdd.n168 0.0180786
R17598 iovdd.n166 iovdd.n165 0.0180786
R17599 iovdd.n165 iovdd.n114 0.0180786
R17600 iovdd.n1356 iovdd.n117 0.0180786
R17601 iovdd.n117 iovdd.n113 0.0180786
R17602 iovdd.n168 iovdd.n166 0.0180786
R17603 iovdd.n1330 iovdd.n164 0.0180786
R17604 iovdd.n171 iovdd.n169 0.0180786
R17605 iovdd.n1331 iovdd.n162 0.0180786
R17606 iovdd.n174 iovdd.n172 0.0180786
R17607 iovdd.n1332 iovdd.n160 0.0180786
R17608 iovdd.n177 iovdd.n175 0.0180786
R17609 iovdd.n1333 iovdd.n158 0.0180786
R17610 iovdd.n180 iovdd.n178 0.0180786
R17611 iovdd.n1334 iovdd.n156 0.0180786
R17612 iovdd.n183 iovdd.n181 0.0180786
R17613 iovdd.n1335 iovdd.n154 0.0180786
R17614 iovdd.n186 iovdd.n184 0.0180786
R17615 iovdd.n1336 iovdd.n152 0.0180786
R17616 iovdd.n189 iovdd.n187 0.0180786
R17617 iovdd.n1337 iovdd.n150 0.0180786
R17618 iovdd.n192 iovdd.n190 0.0180786
R17619 iovdd.n1338 iovdd.n148 0.0180786
R17620 iovdd.n195 iovdd.n193 0.0180786
R17621 iovdd.n1339 iovdd.n146 0.0180786
R17622 iovdd.n198 iovdd.n196 0.0180786
R17623 iovdd.n1340 iovdd.n144 0.0180786
R17624 iovdd.n201 iovdd.n199 0.0180786
R17625 iovdd.n1341 iovdd.n142 0.0180786
R17626 iovdd.n204 iovdd.n202 0.0180786
R17627 iovdd.n1342 iovdd.n140 0.0180786
R17628 iovdd.n207 iovdd.n205 0.0180786
R17629 iovdd.n1343 iovdd.n138 0.0180786
R17630 iovdd.n210 iovdd.n208 0.0180786
R17631 iovdd.n1344 iovdd.n136 0.0180786
R17632 iovdd.n213 iovdd.n211 0.0180786
R17633 iovdd.n1345 iovdd.n134 0.0180786
R17634 iovdd.n216 iovdd.n214 0.0180786
R17635 iovdd.n1346 iovdd.n132 0.0180786
R17636 iovdd.n219 iovdd.n217 0.0180786
R17637 iovdd.n1347 iovdd.n130 0.0180786
R17638 iovdd.n222 iovdd.n220 0.0180786
R17639 iovdd.n1348 iovdd.n128 0.0180786
R17640 iovdd.n225 iovdd.n223 0.0180786
R17641 iovdd.n1349 iovdd.n126 0.0180786
R17642 iovdd.n228 iovdd.n226 0.0180786
R17643 iovdd.n1350 iovdd.n124 0.0180786
R17644 iovdd.n231 iovdd.n229 0.0180786
R17645 iovdd.n1351 iovdd.n122 0.0180786
R17646 iovdd.n234 iovdd.n232 0.0180786
R17647 iovdd.n1352 iovdd.n120 0.0180786
R17648 iovdd.n1354 iovdd.n237 0.0180786
R17649 iovdd.n1356 iovdd.n114 0.0180786
R17650 iovdd.n1300 iovdd.n401 0.0180786
R17651 iovdd.n1298 iovdd.n400 0.0180786
R17652 iovdd.n1281 iovdd.n404 0.0180786
R17653 iovdd.n402 iovdd.n398 0.0180786
R17654 iovdd.n1280 iovdd.n407 0.0180786
R17655 iovdd.n405 iovdd.n396 0.0180786
R17656 iovdd.n1279 iovdd.n410 0.0180786
R17657 iovdd.n408 iovdd.n394 0.0180786
R17658 iovdd.n1303 iovdd.n1302 0.0180786
R17659 iovdd.n411 iovdd.n392 0.0180786
R17660 iovdd.n1305 iovdd.n390 0.0180786
R17661 iovdd.n1251 iovdd.n1249 0.0180786
R17662 iovdd.n1248 iovdd.n560 0.0180786
R17663 iovdd.n1254 iovdd.n1252 0.0180786
R17664 iovdd.n1246 iovdd.n561 0.0180786
R17665 iovdd.n1257 iovdd.n1255 0.0180786
R17666 iovdd.n1244 iovdd.n562 0.0180786
R17667 iovdd.n1260 iovdd.n1258 0.0180786
R17668 iovdd.n1242 iovdd.n563 0.0180786
R17669 iovdd.n1262 iovdd.n566 0.0180786
R17670 iovdd.n1263 iovdd.n565 0.0180786
R17671 iovdd.n564 iovdd.n388 0.0180786
R17672 iovdd.n786 iovdd.n785 0.0180786
R17673 iovdd.n784 iovdd.n775 0.0180786
R17674 iovdd.n788 iovdd.n787 0.0180786
R17675 iovdd.n783 iovdd.n776 0.0180786
R17676 iovdd.n1232 iovdd.n789 0.0180786
R17677 iovdd.n782 iovdd.n777 0.0180786
R17678 iovdd.n1234 iovdd.n779 0.0180786
R17679 iovdd.n1235 iovdd.n778 0.0180786
R17680 iovdd.n1237 iovdd.n569 0.0180786
R17681 iovdd.n773 iovdd.n568 0.0180786
R17682 iovdd.n770 iovdd.n387 0.0180786
R17683 iovdd.n399 iovdd.n56 0.0179603
R17684 iovdd.n227 iovdd.n69 0.0179603
R17685 iovdd.n197 iovdd.n90 0.0179603
R17686 iovdd.n176 iovdd.n103 0.0179603
R17687 iovdd.n1247 iovdd.n354 0.0179603
R17688 iovdd.n539 iovdd.n341 0.0179603
R17689 iovdd.n509 iovdd.n320 0.0179603
R17690 iovdd.n488 iovdd.n307 0.0179603
R17691 iovdd.n849 iovdd.n848 0.0179603
R17692 iovdd.n1175 iovdd.n833 0.0179603
R17693 iovdd.n1155 iovdd.n812 0.0179603
R17694 iovdd.n1141 iovdd.n799 0.0179603
R17695 iovdd.n1289 iovdd.n61 0.0175485
R17696 iovdd.n238 iovdd.n64 0.0175485
R17697 iovdd.n188 iovdd.n95 0.0175485
R17698 iovdd.n185 iovdd.n98 0.0175485
R17699 iovdd.n429 iovdd.n349 0.0175485
R17700 iovdd.n549 iovdd.n346 0.0175485
R17701 iovdd.n500 iovdd.n315 0.0175485
R17702 iovdd.n497 iovdd.n312 0.0175485
R17703 iovdd.n1191 iovdd.n841 0.0175485
R17704 iovdd.n1219 iovdd.n838 0.0175485
R17705 iovdd.n1149 iovdd.n807 0.0175485
R17706 iovdd.n1147 iovdd.n804 0.0175485
R17707 iovdd.n1311 iovdd.n296 0.0175485
R17708 iovdd.n133 iovdd.n78 0.0170873
R17709 iovdd.n135 iovdd.n81 0.0170873
R17710 iovdd.n447 iovdd.n332 0.0170873
R17711 iovdd.n449 iovdd.n329 0.0170873
R17712 iovdd.n1105 iovdd.n824 0.0170873
R17713 iovdd.n1107 iovdd.n821 0.0170873
R17714 iovdd.n403 iovdd.n55 0.0166755
R17715 iovdd.n125 iovdd.n70 0.0166755
R17716 iovdd.n143 iovdd.n89 0.0166755
R17717 iovdd.n159 iovdd.n104 0.0166755
R17718 iovdd.n1253 iovdd.n355 0.0166755
R17719 iovdd.n439 iovdd.n340 0.0166755
R17720 iovdd.n457 iovdd.n321 0.0166755
R17721 iovdd.n473 iovdd.n306 0.0166755
R17722 iovdd.n851 iovdd.n850 0.0166755
R17723 iovdd.n1097 iovdd.n832 0.0166755
R17724 iovdd.n1115 iovdd.n813 0.0166755
R17725 iovdd.n1131 iovdd.n798 0.0166755
R17726 iovdd.n397 iovdd.n53 0.0162143
R17727 iovdd.n224 iovdd.n72 0.0162143
R17728 iovdd.n200 iovdd.n87 0.0162143
R17729 iovdd.n173 iovdd.n106 0.0162143
R17730 iovdd.n1245 iovdd.n357 0.0162143
R17731 iovdd.n536 iovdd.n338 0.0162143
R17732 iovdd.n512 iovdd.n323 0.0162143
R17733 iovdd.n485 iovdd.n304 0.0162143
R17734 iovdd.n1230 iovdd.n791 0.0162143
R17735 iovdd.n1173 iovdd.n830 0.0162143
R17736 iovdd.n1157 iovdd.n815 0.0162143
R17737 iovdd.n1139 iovdd.n796 0.0162143
R17738 iovdd.n524 iovdd.n331 0.0158025
R17739 iovdd.n1165 iovdd.n822 0.0158025
R17740 iovdd.n212 iovdd.n79 0.0158025
R17741 iovdd.n235 iovdd.n62 0.0153413
R17742 iovdd.n235 iovdd.n63 0.0153413
R17743 iovdd.n151 iovdd.n96 0.0153413
R17744 iovdd.n151 iovdd.n97 0.0153413
R17745 iovdd.n432 iovdd.n348 0.0153413
R17746 iovdd.n432 iovdd.n347 0.0153413
R17747 iovdd.n465 iovdd.n314 0.0153413
R17748 iovdd.n465 iovdd.n313 0.0153413
R17749 iovdd.n1193 iovdd.n840 0.0153413
R17750 iovdd.n1193 iovdd.n839 0.0153413
R17751 iovdd.n1123 iovdd.n806 0.0153413
R17752 iovdd.n1123 iovdd.n805 0.0153413
R17753 iovdd.n1310 iovdd.n275 0.0153413
R17754 iovdd.n277 iovdd.n275 0.0153413
R17755 iovdd.n397 iovdd.n54 0.0144683
R17756 iovdd.n224 iovdd.n71 0.0144683
R17757 iovdd.n200 iovdd.n88 0.0144683
R17758 iovdd.n173 iovdd.n105 0.0144683
R17759 iovdd.n1245 iovdd.n356 0.0144683
R17760 iovdd.n536 iovdd.n339 0.0144683
R17761 iovdd.n512 iovdd.n322 0.0144683
R17762 iovdd.n485 iovdd.n305 0.0144683
R17763 iovdd.n852 iovdd.n791 0.0144683
R17764 iovdd.n1173 iovdd.n831 0.0144683
R17765 iovdd.n1157 iovdd.n814 0.0144683
R17766 iovdd.n1139 iovdd.n797 0.0144683
R17767 iovdd.n135 iovdd.n80 0.0135952
R17768 iovdd.n449 iovdd.n330 0.0135952
R17769 iovdd.n1105 iovdd.n823 0.0135952
R17770 iovdd.n116 iovdd 0.0127222
R17771 iovdd.n289 iovdd 0.0109762
R17772 iovdd.n1225 iovdd.n0 0.00923016
R17773 iovdd.n1228 iovdd.n1227 0.00835714
R17774 iovdd.n1357 iovdd.n45 0.00835714
R17775 iovdd.n1239 iovdd.n412 0.00748413
R17776 iovdd.n1357 iovdd.n112 0.00748413
R17777 iovdd.n1240 iovdd.n1239 0.00748413
R17778 iovdd.n298 iovdd.n275 0.00748413
R17779 iovdd.n1239 iovdd.n1238 0.00748413
R17780 iovdd.n1227 iovdd.n859 0.00748413
R17781 iovdd.n943 iovdd.n936 0.00740196
R17782 iovdd.n947 iovdd.n936 0.00740196
R17783 iovdd.n947 iovdd.n929 0.00740196
R17784 iovdd.n958 iovdd.n929 0.00740196
R17785 iovdd.n958 iovdd.n927 0.00740196
R17786 iovdd.n962 iovdd.n927 0.00740196
R17787 iovdd.n962 iovdd.n920 0.00740196
R17788 iovdd.n973 iovdd.n920 0.00740196
R17789 iovdd.n973 iovdd.n918 0.00740196
R17790 iovdd.n977 iovdd.n918 0.00740196
R17791 iovdd.n977 iovdd.n911 0.00740196
R17792 iovdd.n988 iovdd.n911 0.00740196
R17793 iovdd.n988 iovdd.n909 0.00740196
R17794 iovdd.n992 iovdd.n909 0.00740196
R17795 iovdd.n992 iovdd.n902 0.00740196
R17796 iovdd.n1003 iovdd.n902 0.00740196
R17797 iovdd.n1003 iovdd.n900 0.00740196
R17798 iovdd.n1007 iovdd.n900 0.00740196
R17799 iovdd.n1007 iovdd.n893 0.00740196
R17800 iovdd.n1018 iovdd.n893 0.00740196
R17801 iovdd.n1018 iovdd.n891 0.00740196
R17802 iovdd.n1022 iovdd.n891 0.00740196
R17803 iovdd.n1022 iovdd.n884 0.00740196
R17804 iovdd.n1033 iovdd.n884 0.00740196
R17805 iovdd.n1033 iovdd.n882 0.00740196
R17806 iovdd.n1037 iovdd.n882 0.00740196
R17807 iovdd.n1037 iovdd.n875 0.00740196
R17808 iovdd.n1048 iovdd.n875 0.00740196
R17809 iovdd.n1048 iovdd.n873 0.00740196
R17810 iovdd.n1052 iovdd.n873 0.00740196
R17811 iovdd.n1052 iovdd.n866 0.00740196
R17812 iovdd.n1063 iovdd.n866 0.00740196
R17813 iovdd.n1063 iovdd.n246 0.00740196
R17814 iovdd.n1315 iovdd.n246 0.00740196
R17815 iovdd.n1315 iovdd.n240 0.00740196
R17816 iovdd.n1327 iovdd.n240 0.00740196
R17817 iovdd.n1327 iovdd.n1326 0.00740196
R17818 iovdd.n946 iovdd.n945 0.00740196
R17819 iovdd.n946 iovdd.n928 0.00740196
R17820 iovdd.n959 iovdd.n928 0.00740196
R17821 iovdd.n960 iovdd.n959 0.00740196
R17822 iovdd.n961 iovdd.n960 0.00740196
R17823 iovdd.n961 iovdd.n919 0.00740196
R17824 iovdd.n974 iovdd.n919 0.00740196
R17825 iovdd.n975 iovdd.n974 0.00740196
R17826 iovdd.n976 iovdd.n975 0.00740196
R17827 iovdd.n976 iovdd.n910 0.00740196
R17828 iovdd.n989 iovdd.n910 0.00740196
R17829 iovdd.n990 iovdd.n989 0.00740196
R17830 iovdd.n991 iovdd.n990 0.00740196
R17831 iovdd.n991 iovdd.n901 0.00740196
R17832 iovdd.n1004 iovdd.n901 0.00740196
R17833 iovdd.n1005 iovdd.n1004 0.00740196
R17834 iovdd.n1006 iovdd.n1005 0.00740196
R17835 iovdd.n1006 iovdd.n892 0.00740196
R17836 iovdd.n1019 iovdd.n892 0.00740196
R17837 iovdd.n1020 iovdd.n1019 0.00740196
R17838 iovdd.n1021 iovdd.n1020 0.00740196
R17839 iovdd.n1021 iovdd.n883 0.00740196
R17840 iovdd.n1034 iovdd.n883 0.00740196
R17841 iovdd.n1035 iovdd.n1034 0.00740196
R17842 iovdd.n1036 iovdd.n1035 0.00740196
R17843 iovdd.n1036 iovdd.n874 0.00740196
R17844 iovdd.n1049 iovdd.n874 0.00740196
R17845 iovdd.n1050 iovdd.n1049 0.00740196
R17846 iovdd.n1051 iovdd.n1050 0.00740196
R17847 iovdd.n1051 iovdd.n865 0.00740196
R17848 iovdd.n1064 iovdd.n865 0.00740196
R17849 iovdd.n1314 iovdd.n247 0.00740196
R17850 iovdd.n1328 iovdd.n239 0.00740196
R17851 iovdd.n651 iovdd.n650 0.00740196
R17852 iovdd.n651 iovdd.n633 0.00740196
R17853 iovdd.n664 iovdd.n633 0.00740196
R17854 iovdd.n665 iovdd.n664 0.00740196
R17855 iovdd.n666 iovdd.n665 0.00740196
R17856 iovdd.n666 iovdd.n624 0.00740196
R17857 iovdd.n679 iovdd.n624 0.00740196
R17858 iovdd.n680 iovdd.n679 0.00740196
R17859 iovdd.n681 iovdd.n680 0.00740196
R17860 iovdd.n681 iovdd.n615 0.00740196
R17861 iovdd.n694 iovdd.n615 0.00740196
R17862 iovdd.n695 iovdd.n694 0.00740196
R17863 iovdd.n696 iovdd.n695 0.00740196
R17864 iovdd.n696 iovdd.n606 0.00740196
R17865 iovdd.n709 iovdd.n606 0.00740196
R17866 iovdd.n710 iovdd.n709 0.00740196
R17867 iovdd.n711 iovdd.n710 0.00740196
R17868 iovdd.n711 iovdd.n597 0.00740196
R17869 iovdd.n724 iovdd.n597 0.00740196
R17870 iovdd.n725 iovdd.n724 0.00740196
R17871 iovdd.n726 iovdd.n725 0.00740196
R17872 iovdd.n726 iovdd.n588 0.00740196
R17873 iovdd.n739 iovdd.n588 0.00740196
R17874 iovdd.n740 iovdd.n739 0.00740196
R17875 iovdd.n741 iovdd.n740 0.00740196
R17876 iovdd.n741 iovdd.n579 0.00740196
R17877 iovdd.n754 iovdd.n579 0.00740196
R17878 iovdd.n755 iovdd.n754 0.00740196
R17879 iovdd.n756 iovdd.n755 0.00740196
R17880 iovdd.n756 iovdd.n570 0.00740196
R17881 iovdd.n769 iovdd.n570 0.00740196
R17882 iovdd.n1265 iovdd.n422 0.00740196
R17883 iovdd.n1278 iovdd.n413 0.00740196
R17884 iovdd.n648 iovdd.n641 0.00740196
R17885 iovdd.n652 iovdd.n641 0.00740196
R17886 iovdd.n652 iovdd.n634 0.00740196
R17887 iovdd.n663 iovdd.n634 0.00740196
R17888 iovdd.n663 iovdd.n632 0.00740196
R17889 iovdd.n667 iovdd.n632 0.00740196
R17890 iovdd.n667 iovdd.n625 0.00740196
R17891 iovdd.n678 iovdd.n625 0.00740196
R17892 iovdd.n678 iovdd.n623 0.00740196
R17893 iovdd.n682 iovdd.n623 0.00740196
R17894 iovdd.n682 iovdd.n616 0.00740196
R17895 iovdd.n693 iovdd.n616 0.00740196
R17896 iovdd.n693 iovdd.n614 0.00740196
R17897 iovdd.n697 iovdd.n614 0.00740196
R17898 iovdd.n697 iovdd.n607 0.00740196
R17899 iovdd.n708 iovdd.n607 0.00740196
R17900 iovdd.n708 iovdd.n605 0.00740196
R17901 iovdd.n712 iovdd.n605 0.00740196
R17902 iovdd.n712 iovdd.n598 0.00740196
R17903 iovdd.n723 iovdd.n598 0.00740196
R17904 iovdd.n723 iovdd.n596 0.00740196
R17905 iovdd.n727 iovdd.n596 0.00740196
R17906 iovdd.n727 iovdd.n589 0.00740196
R17907 iovdd.n738 iovdd.n589 0.00740196
R17908 iovdd.n738 iovdd.n587 0.00740196
R17909 iovdd.n742 iovdd.n587 0.00740196
R17910 iovdd.n742 iovdd.n580 0.00740196
R17911 iovdd.n753 iovdd.n580 0.00740196
R17912 iovdd.n753 iovdd.n578 0.00740196
R17913 iovdd.n757 iovdd.n578 0.00740196
R17914 iovdd.n757 iovdd.n571 0.00740196
R17915 iovdd.n768 iovdd.n571 0.00740196
R17916 iovdd.n768 iovdd.n421 0.00740196
R17917 iovdd.n1266 iovdd.n421 0.00740196
R17918 iovdd.n1266 iovdd.n414 0.00740196
R17919 iovdd.n1277 iovdd.n414 0.00740196
R17920 iovdd.n1277 iovdd.n415 0.00740196
R17921 iovdd.n1355 iovdd 0.00671176
R17922 iovdd.n863 iovdd.n858 0.0057381
R17923 iovdd.n116 iovdd.n44 0.0057381
R17924 iovdd.n1353 iovdd.n1328 0.0047102
R17925 iovdd.n1301 iovdd.n1278 0.0047102
R17926 iovdd.n944 iovdd.n943 0.00442211
R17927 iovdd.n649 iovdd.n648 0.00442211
R17928 iovdd iovdd.n0 0.00399206
R17929 iovdd.n942 iovdd.n937 0.00395098
R17930 iovdd.n942 iovdd.n941 0.00395098
R17931 iovdd.n941 iovdd.n938 0.00395098
R17932 iovdd.n938 iovdd.n935 0.00395098
R17933 iovdd.n948 iovdd.n935 0.00395098
R17934 iovdd.n950 iovdd.n948 0.00395098
R17935 iovdd.n950 iovdd.n949 0.00395098
R17936 iovdd.n949 iovdd.n930 0.00395098
R17937 iovdd.n957 iovdd.n930 0.00395098
R17938 iovdd.n957 iovdd.n956 0.00395098
R17939 iovdd.n956 iovdd.n931 0.00395098
R17940 iovdd.n931 iovdd.n926 0.00395098
R17941 iovdd.n963 iovdd.n926 0.00395098
R17942 iovdd.n965 iovdd.n963 0.00395098
R17943 iovdd.n965 iovdd.n964 0.00395098
R17944 iovdd.n964 iovdd.n921 0.00395098
R17945 iovdd.n972 iovdd.n921 0.00395098
R17946 iovdd.n972 iovdd.n971 0.00395098
R17947 iovdd.n971 iovdd.n922 0.00395098
R17948 iovdd.n922 iovdd.n917 0.00395098
R17949 iovdd.n978 iovdd.n917 0.00395098
R17950 iovdd.n980 iovdd.n978 0.00395098
R17951 iovdd.n980 iovdd.n979 0.00395098
R17952 iovdd.n979 iovdd.n912 0.00395098
R17953 iovdd.n987 iovdd.n912 0.00395098
R17954 iovdd.n987 iovdd.n986 0.00395098
R17955 iovdd.n986 iovdd.n913 0.00395098
R17956 iovdd.n913 iovdd.n908 0.00395098
R17957 iovdd.n993 iovdd.n908 0.00395098
R17958 iovdd.n995 iovdd.n993 0.00395098
R17959 iovdd.n995 iovdd.n994 0.00395098
R17960 iovdd.n994 iovdd.n903 0.00395098
R17961 iovdd.n1002 iovdd.n903 0.00395098
R17962 iovdd.n1002 iovdd.n1001 0.00395098
R17963 iovdd.n1001 iovdd.n904 0.00395098
R17964 iovdd.n904 iovdd.n899 0.00395098
R17965 iovdd.n1008 iovdd.n899 0.00395098
R17966 iovdd.n1010 iovdd.n1008 0.00395098
R17967 iovdd.n1010 iovdd.n1009 0.00395098
R17968 iovdd.n1009 iovdd.n894 0.00395098
R17969 iovdd.n1017 iovdd.n894 0.00395098
R17970 iovdd.n1017 iovdd.n1016 0.00395098
R17971 iovdd.n1016 iovdd.n895 0.00395098
R17972 iovdd.n895 iovdd.n890 0.00395098
R17973 iovdd.n1023 iovdd.n890 0.00395098
R17974 iovdd.n1025 iovdd.n1023 0.00395098
R17975 iovdd.n1025 iovdd.n1024 0.00395098
R17976 iovdd.n1024 iovdd.n885 0.00395098
R17977 iovdd.n1032 iovdd.n885 0.00395098
R17978 iovdd.n1032 iovdd.n1031 0.00395098
R17979 iovdd.n1031 iovdd.n886 0.00395098
R17980 iovdd.n886 iovdd.n881 0.00395098
R17981 iovdd.n1038 iovdd.n881 0.00395098
R17982 iovdd.n1040 iovdd.n1038 0.00395098
R17983 iovdd.n1040 iovdd.n1039 0.00395098
R17984 iovdd.n1039 iovdd.n876 0.00395098
R17985 iovdd.n1047 iovdd.n876 0.00395098
R17986 iovdd.n1047 iovdd.n1046 0.00395098
R17987 iovdd.n1046 iovdd.n877 0.00395098
R17988 iovdd.n877 iovdd.n872 0.00395098
R17989 iovdd.n1053 iovdd.n872 0.00395098
R17990 iovdd.n1055 iovdd.n1053 0.00395098
R17991 iovdd.n1055 iovdd.n1054 0.00395098
R17992 iovdd.n1054 iovdd.n867 0.00395098
R17993 iovdd.n1062 iovdd.n867 0.00395098
R17994 iovdd.n1062 iovdd.n1061 0.00395098
R17995 iovdd.n1061 iovdd.n868 0.00395098
R17996 iovdd.n868 iovdd.n245 0.00395098
R17997 iovdd.n1316 iovdd.n245 0.00395098
R17998 iovdd.n1319 iovdd.n1316 0.00395098
R17999 iovdd.n1319 iovdd.n1318 0.00395098
R18000 iovdd.n1318 iovdd.n1317 0.00395098
R18001 iovdd.n1317 iovdd.n241 0.00395098
R18002 iovdd.n1325 iovdd.n241 0.00395098
R18003 iovdd.n647 iovdd.n642 0.00395098
R18004 iovdd.n647 iovdd.n646 0.00395098
R18005 iovdd.n646 iovdd.n643 0.00395098
R18006 iovdd.n643 iovdd.n640 0.00395098
R18007 iovdd.n653 iovdd.n640 0.00395098
R18008 iovdd.n655 iovdd.n653 0.00395098
R18009 iovdd.n655 iovdd.n654 0.00395098
R18010 iovdd.n654 iovdd.n635 0.00395098
R18011 iovdd.n662 iovdd.n635 0.00395098
R18012 iovdd.n662 iovdd.n661 0.00395098
R18013 iovdd.n661 iovdd.n636 0.00395098
R18014 iovdd.n636 iovdd.n631 0.00395098
R18015 iovdd.n668 iovdd.n631 0.00395098
R18016 iovdd.n670 iovdd.n668 0.00395098
R18017 iovdd.n670 iovdd.n669 0.00395098
R18018 iovdd.n669 iovdd.n626 0.00395098
R18019 iovdd.n677 iovdd.n626 0.00395098
R18020 iovdd.n677 iovdd.n676 0.00395098
R18021 iovdd.n676 iovdd.n627 0.00395098
R18022 iovdd.n627 iovdd.n622 0.00395098
R18023 iovdd.n683 iovdd.n622 0.00395098
R18024 iovdd.n685 iovdd.n683 0.00395098
R18025 iovdd.n685 iovdd.n684 0.00395098
R18026 iovdd.n684 iovdd.n617 0.00395098
R18027 iovdd.n692 iovdd.n617 0.00395098
R18028 iovdd.n692 iovdd.n691 0.00395098
R18029 iovdd.n691 iovdd.n618 0.00395098
R18030 iovdd.n618 iovdd.n613 0.00395098
R18031 iovdd.n698 iovdd.n613 0.00395098
R18032 iovdd.n700 iovdd.n698 0.00395098
R18033 iovdd.n700 iovdd.n699 0.00395098
R18034 iovdd.n699 iovdd.n608 0.00395098
R18035 iovdd.n707 iovdd.n608 0.00395098
R18036 iovdd.n707 iovdd.n706 0.00395098
R18037 iovdd.n706 iovdd.n609 0.00395098
R18038 iovdd.n609 iovdd.n604 0.00395098
R18039 iovdd.n713 iovdd.n604 0.00395098
R18040 iovdd.n715 iovdd.n713 0.00395098
R18041 iovdd.n715 iovdd.n714 0.00395098
R18042 iovdd.n714 iovdd.n599 0.00395098
R18043 iovdd.n722 iovdd.n599 0.00395098
R18044 iovdd.n722 iovdd.n721 0.00395098
R18045 iovdd.n721 iovdd.n600 0.00395098
R18046 iovdd.n600 iovdd.n595 0.00395098
R18047 iovdd.n728 iovdd.n595 0.00395098
R18048 iovdd.n730 iovdd.n728 0.00395098
R18049 iovdd.n730 iovdd.n729 0.00395098
R18050 iovdd.n729 iovdd.n590 0.00395098
R18051 iovdd.n737 iovdd.n590 0.00395098
R18052 iovdd.n737 iovdd.n736 0.00395098
R18053 iovdd.n736 iovdd.n591 0.00395098
R18054 iovdd.n591 iovdd.n586 0.00395098
R18055 iovdd.n743 iovdd.n586 0.00395098
R18056 iovdd.n745 iovdd.n743 0.00395098
R18057 iovdd.n745 iovdd.n744 0.00395098
R18058 iovdd.n744 iovdd.n581 0.00395098
R18059 iovdd.n752 iovdd.n581 0.00395098
R18060 iovdd.n752 iovdd.n751 0.00395098
R18061 iovdd.n751 iovdd.n582 0.00395098
R18062 iovdd.n582 iovdd.n577 0.00395098
R18063 iovdd.n758 iovdd.n577 0.00395098
R18064 iovdd.n760 iovdd.n758 0.00395098
R18065 iovdd.n760 iovdd.n759 0.00395098
R18066 iovdd.n759 iovdd.n572 0.00395098
R18067 iovdd.n767 iovdd.n572 0.00395098
R18068 iovdd.n767 iovdd.n766 0.00395098
R18069 iovdd.n766 iovdd.n573 0.00395098
R18070 iovdd.n573 iovdd.n420 0.00395098
R18071 iovdd.n1267 iovdd.n420 0.00395098
R18072 iovdd.n1269 iovdd.n1267 0.00395098
R18073 iovdd.n1269 iovdd.n1268 0.00395098
R18074 iovdd.n1268 iovdd.n416 0.00395098
R18075 iovdd.n1276 iovdd.n416 0.00395098
R18076 iovdd.n1276 iovdd.n1275 0.00395098
R18077 iovdd.n1239 iovdd.n49 0.00360916
R18078 iovdd.n1306 iovdd.n375 0.00339474
R18079 iovdd.n1218 iovdd.n247 0.00326078
R18080 iovdd.n1233 iovdd.n422 0.00326078
R18081 iovdd.n1314 iovdd.n1313 0.00298471
R18082 iovdd.n1265 iovdd.n1264 0.00298471
R18083 iovdd.n772 iovdd.n375 0.00285867
R18084 iovdd.n1274 iovdd 0.00261765
R18085 iovdd.n290 iovdd.n289 0.00224603
R18086 iovdd.n1236 iovdd.n774 0.00219098
R18087 iovdd.n1264 iovdd.n559 0.00219098
R18088 iovdd.n1261 iovdd.n559 0.00219098
R18089 iovdd.n1273 iovdd 0.00196667
R18090 iovdd.n1323 iovdd 0.00196667
R18091 iovdd.n940 iovdd.n934 0.00191176
R18092 iovdd.n951 iovdd.n934 0.00191176
R18093 iovdd.n951 iovdd.n932 0.00191176
R18094 iovdd.n955 iovdd.n932 0.00191176
R18095 iovdd.n955 iovdd.n925 0.00191176
R18096 iovdd.n966 iovdd.n925 0.00191176
R18097 iovdd.n966 iovdd.n923 0.00191176
R18098 iovdd.n970 iovdd.n923 0.00191176
R18099 iovdd.n970 iovdd.n916 0.00191176
R18100 iovdd.n981 iovdd.n916 0.00191176
R18101 iovdd.n981 iovdd.n914 0.00191176
R18102 iovdd.n985 iovdd.n914 0.00191176
R18103 iovdd.n985 iovdd.n907 0.00191176
R18104 iovdd.n996 iovdd.n907 0.00191176
R18105 iovdd.n996 iovdd.n905 0.00191176
R18106 iovdd.n1000 iovdd.n905 0.00191176
R18107 iovdd.n1000 iovdd.n898 0.00191176
R18108 iovdd.n1011 iovdd.n898 0.00191176
R18109 iovdd.n1011 iovdd.n896 0.00191176
R18110 iovdd.n1015 iovdd.n896 0.00191176
R18111 iovdd.n1015 iovdd.n889 0.00191176
R18112 iovdd.n1026 iovdd.n889 0.00191176
R18113 iovdd.n1026 iovdd.n887 0.00191176
R18114 iovdd.n1030 iovdd.n887 0.00191176
R18115 iovdd.n1030 iovdd.n880 0.00191176
R18116 iovdd.n1041 iovdd.n880 0.00191176
R18117 iovdd.n1041 iovdd.n878 0.00191176
R18118 iovdd.n1045 iovdd.n878 0.00191176
R18119 iovdd.n1045 iovdd.n871 0.00191176
R18120 iovdd.n1056 iovdd.n871 0.00191176
R18121 iovdd.n1056 iovdd.n869 0.00191176
R18122 iovdd.n1060 iovdd.n869 0.00191176
R18123 iovdd.n1060 iovdd.n244 0.00191176
R18124 iovdd.n1320 iovdd.n244 0.00191176
R18125 iovdd.n1320 iovdd.n242 0.00191176
R18126 iovdd.n1324 iovdd.n242 0.00191176
R18127 iovdd.n645 iovdd.n639 0.00191176
R18128 iovdd.n656 iovdd.n639 0.00191176
R18129 iovdd.n656 iovdd.n637 0.00191176
R18130 iovdd.n660 iovdd.n637 0.00191176
R18131 iovdd.n660 iovdd.n630 0.00191176
R18132 iovdd.n671 iovdd.n630 0.00191176
R18133 iovdd.n671 iovdd.n628 0.00191176
R18134 iovdd.n675 iovdd.n628 0.00191176
R18135 iovdd.n675 iovdd.n621 0.00191176
R18136 iovdd.n686 iovdd.n621 0.00191176
R18137 iovdd.n686 iovdd.n619 0.00191176
R18138 iovdd.n690 iovdd.n619 0.00191176
R18139 iovdd.n690 iovdd.n612 0.00191176
R18140 iovdd.n701 iovdd.n612 0.00191176
R18141 iovdd.n701 iovdd.n610 0.00191176
R18142 iovdd.n705 iovdd.n610 0.00191176
R18143 iovdd.n705 iovdd.n603 0.00191176
R18144 iovdd.n716 iovdd.n603 0.00191176
R18145 iovdd.n716 iovdd.n601 0.00191176
R18146 iovdd.n720 iovdd.n601 0.00191176
R18147 iovdd.n720 iovdd.n594 0.00191176
R18148 iovdd.n731 iovdd.n594 0.00191176
R18149 iovdd.n731 iovdd.n592 0.00191176
R18150 iovdd.n735 iovdd.n592 0.00191176
R18151 iovdd.n735 iovdd.n585 0.00191176
R18152 iovdd.n746 iovdd.n585 0.00191176
R18153 iovdd.n746 iovdd.n583 0.00191176
R18154 iovdd.n750 iovdd.n583 0.00191176
R18155 iovdd.n750 iovdd.n576 0.00191176
R18156 iovdd.n761 iovdd.n576 0.00191176
R18157 iovdd.n761 iovdd.n574 0.00191176
R18158 iovdd.n765 iovdd.n574 0.00191176
R18159 iovdd.n765 iovdd.n419 0.00191176
R18160 iovdd.n1270 iovdd.n419 0.00191176
R18161 iovdd.n1270 iovdd.n417 0.00191176
R18162 iovdd.n1274 iovdd.n417 0.00191176
R18163 iovdd.n1294 iovdd.n389 0.00189683
R18164 iovdd.n1286 iovdd.n115 0.00189683
R18165 iovdd.n1183 iovdd.n774 0.00189683
R18166 iovdd.n1221 iovdd.n1090 0.00189683
R18167 iovdd.n559 iovdd.n558 0.00189683
R18168 iovdd.n552 iovdd.n431 0.00189683
R18169 iovdd.n1222 iovdd.n1221 0.00184541
R18170 iovdd.n1218 iovdd.n864 0.00184541
R18171 iovdd.n431 iovdd.n248 0.00184541
R18172 iovdd.n548 iovdd.n431 0.00184541
R18173 iovdd.n1329 iovdd.n115 0.00184541
R18174 iovdd.n548 iovdd.n547 0.00184541
R18175 iovdd.n1313 iovdd.n248 0.00184541
R18176 iovdd.n1223 iovdd.n1222 0.00184541
R18177 iovdd.n1221 iovdd.n864 0.00184541
R18178 iovdd.n1353 iovdd.n1329 0.00184541
R18179 iovdd.n1233 iovdd.n781 0.00184541
R18180 iovdd.n1297 iovdd.n389 0.00184541
R18181 iovdd.n1301 iovdd.n1297 0.00184541
R18182 iovdd.n781 iovdd.n774 0.00184541
R18183 iovdd.n772 iovdd.n49 0.00178655
R18184 iovdd.n940 iovdd.n939 0.0016983
R18185 iovdd.n645 iovdd.n644 0.0016983
R18186 iovdd.n547 iovdd.n239 0.00153529
R18187 iovdd.n1261 iovdd.n413 0.00153529
R18188 iovdd.n118 iovdd.n115 0.00150078
R18189 iovdd.n391 iovdd.n389 0.00150078
R18190 iovdd.n657 iovdd.n638 0.00147778
R18191 iovdd.n658 iovdd.n657 0.00147778
R18192 iovdd.n659 iovdd.n658 0.00147778
R18193 iovdd.n659 iovdd.n629 0.00147778
R18194 iovdd.n672 iovdd.n629 0.00147778
R18195 iovdd.n673 iovdd.n672 0.00147778
R18196 iovdd.n674 iovdd.n673 0.00147778
R18197 iovdd.n674 iovdd.n620 0.00147778
R18198 iovdd.n687 iovdd.n620 0.00147778
R18199 iovdd.n688 iovdd.n687 0.00147778
R18200 iovdd.n689 iovdd.n688 0.00147778
R18201 iovdd.n689 iovdd.n611 0.00147778
R18202 iovdd.n702 iovdd.n611 0.00147778
R18203 iovdd.n703 iovdd.n702 0.00147778
R18204 iovdd.n704 iovdd.n703 0.00147778
R18205 iovdd.n704 iovdd.n602 0.00147778
R18206 iovdd.n717 iovdd.n602 0.00147778
R18207 iovdd.n718 iovdd.n717 0.00147778
R18208 iovdd.n719 iovdd.n718 0.00147778
R18209 iovdd.n719 iovdd.n593 0.00147778
R18210 iovdd.n732 iovdd.n593 0.00147778
R18211 iovdd.n733 iovdd.n732 0.00147778
R18212 iovdd.n734 iovdd.n733 0.00147778
R18213 iovdd.n734 iovdd.n584 0.00147778
R18214 iovdd.n747 iovdd.n584 0.00147778
R18215 iovdd.n748 iovdd.n747 0.00147778
R18216 iovdd.n749 iovdd.n748 0.00147778
R18217 iovdd.n749 iovdd.n575 0.00147778
R18218 iovdd.n762 iovdd.n575 0.00147778
R18219 iovdd.n763 iovdd.n762 0.00147778
R18220 iovdd.n764 iovdd.n763 0.00147778
R18221 iovdd.n764 iovdd.n418 0.00147778
R18222 iovdd.n1271 iovdd.n418 0.00147778
R18223 iovdd.n1272 iovdd.n1271 0.00147778
R18224 iovdd.n1273 iovdd.n1272 0.00147778
R18225 iovdd.n952 iovdd.n933 0.00147778
R18226 iovdd.n953 iovdd.n952 0.00147778
R18227 iovdd.n954 iovdd.n953 0.00147778
R18228 iovdd.n954 iovdd.n924 0.00147778
R18229 iovdd.n967 iovdd.n924 0.00147778
R18230 iovdd.n968 iovdd.n967 0.00147778
R18231 iovdd.n969 iovdd.n968 0.00147778
R18232 iovdd.n969 iovdd.n915 0.00147778
R18233 iovdd.n982 iovdd.n915 0.00147778
R18234 iovdd.n983 iovdd.n982 0.00147778
R18235 iovdd.n984 iovdd.n983 0.00147778
R18236 iovdd.n984 iovdd.n906 0.00147778
R18237 iovdd.n997 iovdd.n906 0.00147778
R18238 iovdd.n998 iovdd.n997 0.00147778
R18239 iovdd.n999 iovdd.n998 0.00147778
R18240 iovdd.n999 iovdd.n897 0.00147778
R18241 iovdd.n1012 iovdd.n897 0.00147778
R18242 iovdd.n1013 iovdd.n1012 0.00147778
R18243 iovdd.n1014 iovdd.n1013 0.00147778
R18244 iovdd.n1014 iovdd.n888 0.00147778
R18245 iovdd.n1027 iovdd.n888 0.00147778
R18246 iovdd.n1028 iovdd.n1027 0.00147778
R18247 iovdd.n1029 iovdd.n1028 0.00147778
R18248 iovdd.n1029 iovdd.n879 0.00147778
R18249 iovdd.n1042 iovdd.n879 0.00147778
R18250 iovdd.n1043 iovdd.n1042 0.00147778
R18251 iovdd.n1044 iovdd.n1043 0.00147778
R18252 iovdd.n1044 iovdd.n870 0.00147778
R18253 iovdd.n1057 iovdd.n870 0.00147778
R18254 iovdd.n1058 iovdd.n1057 0.00147778
R18255 iovdd.n1059 iovdd.n1058 0.00147778
R18256 iovdd.n1059 iovdd.n243 0.00147778
R18257 iovdd.n1321 iovdd.n243 0.00147778
R18258 iovdd.n1322 iovdd.n1321 0.00147778
R18259 iovdd.n1323 iovdd.n1322 0.00147778
R18260 iovdd.n1223 iovdd.n1064 0.00125922
R18261 iovdd.n1236 iovdd.n769 0.00125922
R18262 iovdd.n1307 iovdd.n1306 0.00125049
R18263 iovdd.n1355 iovdd.n118 0.0011902
R18264 iovdd.n1304 iovdd.n391 0.0011902
R18265 iovdd.n1360 iovdd.n1359 0.00101087
R18266 iovdd.n1309 iovdd.n25 0.001
R18267 iovdd.n1229 iovdd.n8 0.001
R18268 iovdd.n363 iovdd.n7 0.001
R18269 iovdd.n376 iovdd.n7 0.001
R18270 iovdd.n857 iovdd.n9 0.001
R18271 iovdd.n377 iovdd.n9 0.001
R18272 iovdd.n364 iovdd.n11 0.001
R18273 iovdd.n378 iovdd.n11 0.001
R18274 iovdd.n365 iovdd.n13 0.001
R18275 iovdd.n379 iovdd.n13 0.001
R18276 iovdd.n366 iovdd.n17 0.001
R18277 iovdd.n380 iovdd.n17 0.001
R18278 iovdd.n367 iovdd.n20 0.001
R18279 iovdd.n381 iovdd.n20 0.001
R18280 iovdd.n368 iovdd.n23 0.001
R18281 iovdd.n1308 iovdd.n23 0.001
R18282 iovdd.n1309 iovdd.n362 0.001
R18283 iovdd.n369 iovdd.n28 0.001
R18284 iovdd.n382 iovdd.n28 0.001
R18285 iovdd.n370 iovdd.n31 0.001
R18286 iovdd.n383 iovdd.n31 0.001
R18287 iovdd.n371 iovdd.n34 0.001
R18288 iovdd.n384 iovdd.n34 0.001
R18289 iovdd.n372 iovdd.n37 0.001
R18290 iovdd.n385 iovdd.n37 0.001
R18291 iovdd.n373 iovdd.n40 0.001
R18292 iovdd.n386 iovdd.n40 0.001
R18293 iovdd.n1359 iovdd.n48 0.001
R18294 iovdd.n1359 iovdd.n47 0.001
R18295 iovdd.n374 iovdd.n43 0.001
R18296 iovdd.n47 iovdd.n4 0.001
R18297 iovdd.n386 iovdd.n42 0.001
R18298 iovdd.n385 iovdd.n39 0.001
R18299 iovdd.n384 iovdd.n36 0.001
R18300 iovdd.n383 iovdd.n33 0.001
R18301 iovdd.n382 iovdd.n30 0.001
R18302 iovdd.n362 iovdd.n27 0.001
R18303 iovdd.n1309 iovdd.n1308 0.001
R18304 iovdd.n381 iovdd.n22 0.001
R18305 iovdd.n380 iovdd.n19 0.001
R18306 iovdd.n379 iovdd.n16 0.001
R18307 iovdd.n378 iovdd.n12 0.001
R18308 iovdd.n377 iovdd.n10 0.001
R18309 iovdd.n1229 iovdd.n376 0.001
R18310 iovdd.n374 iovdd.n4 0.001
R18311 iovdd.n48 iovdd.n42 0.001
R18312 iovdd.n373 iovdd.n39 0.001
R18313 iovdd.n372 iovdd.n36 0.001
R18314 iovdd.n371 iovdd.n33 0.001
R18315 iovdd.n370 iovdd.n30 0.001
R18316 iovdd.n369 iovdd.n27 0.001
R18317 iovdd.n368 iovdd.n22 0.001
R18318 iovdd.n367 iovdd.n19 0.001
R18319 iovdd.n366 iovdd.n16 0.001
R18320 iovdd.n365 iovdd.n12 0.001
R18321 iovdd.n364 iovdd.n10 0.001
R18322 iovdd.n1229 iovdd.n857 0.001
R18323 iovdd.n363 iovdd.n5 0.001
R18324 iovdd.n8 iovdd.n3 0.001
R18325 iovdd.n1361 iovdd.n3 0.001
R18326 iovdd.n1362 iovdd.n2 0.001
R18327 iovdd.n15 iovdd.n14 0.001
R18328 iovdd.n293 iovdd.n18 0.001
R18329 iovdd.n292 iovdd.n21 0.001
R18330 iovdd.n291 iovdd.n24 0.001
R18331 iovdd.n288 iovdd.n25 0.001
R18332 iovdd.n288 iovdd.n26 0.001
R18333 iovdd.n286 iovdd.n29 0.001
R18334 iovdd.n284 iovdd.n32 0.001
R18335 iovdd.n282 iovdd.n35 0.001
R18336 iovdd.n280 iovdd.n38 0.001
R18337 iovdd.n278 iovdd.n41 0.001
R18338 iovdd.n1359 iovdd.n41 0.001
R18339 iovdd.n278 iovdd.n38 0.001
R18340 iovdd.n280 iovdd.n35 0.001
R18341 iovdd.n282 iovdd.n32 0.001
R18342 iovdd.n284 iovdd.n29 0.001
R18343 iovdd.n286 iovdd.n26 0.001
R18344 iovdd.n1309 iovdd.n24 0.001
R18345 iovdd.n1229 iovdd.n6 0.001
R18346 iovdd.n291 iovdd.n21 0.001
R18347 iovdd.n292 iovdd.n18 0.001
R18348 iovdd.n293 iovdd.n15 0.001
R18349 iovdd.n14 iovdd.n2 0.001
R18350 iovdd.n1362 iovdd.n1361 0.001
R18351 vdd.n74 vdd.n73 1.50539
R18352 vdd.n1 vdd.n0 1.5005
R18353 vdd.n69 vdd.n68 1.5005
R18354 vdd.n67 vdd.n66 1.5005
R18355 vdd.n5 vdd.n4 1.5005
R18356 vdd.n61 vdd.n60 1.5005
R18357 vdd.n59 vdd.n58 1.5005
R18358 vdd.n9 vdd.n8 1.5005
R18359 vdd.n53 vdd.n52 1.5005
R18360 vdd.n51 vdd.n50 1.5005
R18361 vdd.n13 vdd.n12 1.5005
R18362 vdd.n45 vdd.n44 1.5005
R18363 vdd.n43 vdd.n42 1.5005
R18364 vdd.n17 vdd.n16 1.5005
R18365 vdd.n37 vdd.n36 1.5005
R18366 vdd.n35 vdd.n34 1.5005
R18367 vdd.n21 vdd.n20 1.5005
R18368 vdd.n29 vdd.n28 1.5005
R18369 vdd.n27 vdd.n26 1.5005
R18370 vdd.n75 vdd 0.6957
R18371 vdd.n73 vdd.n72 0.314786
R18372 vdd.n71 vdd.n70 0.314786
R18373 vdd.n3 vdd.n2 0.314786
R18374 vdd.n65 vdd.n64 0.314786
R18375 vdd.n63 vdd.n62 0.314786
R18376 vdd.n7 vdd.n6 0.314786
R18377 vdd.n57 vdd.n56 0.314786
R18378 vdd.n55 vdd.n54 0.314786
R18379 vdd.n11 vdd.n10 0.314786
R18380 vdd.n49 vdd.n48 0.314786
R18381 vdd.n47 vdd.n46 0.314786
R18382 vdd.n15 vdd.n14 0.314786
R18383 vdd.n41 vdd.n40 0.314786
R18384 vdd.n39 vdd.n38 0.314786
R18385 vdd.n19 vdd.n18 0.314786
R18386 vdd.n33 vdd.n32 0.314786
R18387 vdd.n31 vdd.n30 0.314786
R18388 vdd.n23 vdd.n22 0.314786
R18389 vdd.n24 vdd 0.217715
R18390 vdd.n51 vdd 0.195018
R18391 vdd.n25 vdd.n24 0.146103
R18392 vdd.n26 vdd.n25 0.0354467
R18393 vdd.n25 vdd.n22 0.0314255
R18394 vdd.n28 vdd.n27 0.00921287
R18395 vdd.n28 vdd.n20 0.00921287
R18396 vdd.n35 vdd.n20 0.00921287
R18397 vdd.n36 vdd.n35 0.00921287
R18398 vdd.n36 vdd.n16 0.00921287
R18399 vdd.n43 vdd.n16 0.00921287
R18400 vdd.n44 vdd.n43 0.00921287
R18401 vdd.n44 vdd.n12 0.00921287
R18402 vdd.n51 vdd.n12 0.00921287
R18403 vdd.n52 vdd.n51 0.00921287
R18404 vdd.n52 vdd.n8 0.00921287
R18405 vdd.n59 vdd.n8 0.00921287
R18406 vdd.n60 vdd.n59 0.00921287
R18407 vdd.n60 vdd.n4 0.00921287
R18408 vdd.n67 vdd.n4 0.00921287
R18409 vdd.n68 vdd.n67 0.00921287
R18410 vdd.n68 vdd.n0 0.00921287
R18411 vdd.n74 vdd.n0 0.00921287
R18412 vdd.n26 vdd.n23 0.00538889
R18413 vdd.n29 vdd.n23 0.00538889
R18414 vdd.n30 vdd.n29 0.00538889
R18415 vdd.n30 vdd.n21 0.00538889
R18416 vdd.n33 vdd.n21 0.00538889
R18417 vdd.n34 vdd.n33 0.00538889
R18418 vdd.n34 vdd.n19 0.00538889
R18419 vdd.n37 vdd.n19 0.00538889
R18420 vdd.n38 vdd.n37 0.00538889
R18421 vdd.n38 vdd.n17 0.00538889
R18422 vdd.n41 vdd.n17 0.00538889
R18423 vdd.n42 vdd.n41 0.00538889
R18424 vdd.n42 vdd.n15 0.00538889
R18425 vdd.n45 vdd.n15 0.00538889
R18426 vdd.n46 vdd.n45 0.00538889
R18427 vdd.n46 vdd.n13 0.00538889
R18428 vdd.n49 vdd.n13 0.00538889
R18429 vdd.n50 vdd.n49 0.00538889
R18430 vdd.n50 vdd.n11 0.00538889
R18431 vdd.n53 vdd.n11 0.00538889
R18432 vdd.n54 vdd.n53 0.00538889
R18433 vdd.n54 vdd.n9 0.00538889
R18434 vdd.n57 vdd.n9 0.00538889
R18435 vdd.n58 vdd.n57 0.00538889
R18436 vdd.n58 vdd.n7 0.00538889
R18437 vdd.n61 vdd.n7 0.00538889
R18438 vdd.n62 vdd.n61 0.00538889
R18439 vdd.n62 vdd.n5 0.00538889
R18440 vdd.n65 vdd.n5 0.00538889
R18441 vdd.n66 vdd.n65 0.00538889
R18442 vdd.n66 vdd.n3 0.00538889
R18443 vdd.n69 vdd.n3 0.00538889
R18444 vdd.n70 vdd.n69 0.00538889
R18445 vdd.n70 vdd.n1 0.00538889
R18446 vdd.n73 vdd.n1 0.00538889
R18447 vdd.n27 vdd.n24 0.00485644
R18448 vdd.n75 vdd.n74 0.00485644
R18449 vdd vdd.n75 0.00485644
R18450 vdd.n72 vdd 0.0035
R18451 vdd.n31 vdd.n22 0.0025
R18452 vdd.n32 vdd.n31 0.0025
R18453 vdd.n32 vdd.n18 0.0025
R18454 vdd.n39 vdd.n18 0.0025
R18455 vdd.n40 vdd.n39 0.0025
R18456 vdd.n40 vdd.n14 0.0025
R18457 vdd.n47 vdd.n14 0.0025
R18458 vdd.n48 vdd.n47 0.0025
R18459 vdd.n48 vdd.n10 0.0025
R18460 vdd.n55 vdd.n10 0.0025
R18461 vdd.n56 vdd.n55 0.0025
R18462 vdd.n56 vdd.n6 0.0025
R18463 vdd.n63 vdd.n6 0.0025
R18464 vdd.n64 vdd.n63 0.0025
R18465 vdd.n64 vdd.n2 0.0025
R18466 vdd.n71 vdd.n2 0.0025
R18467 vdd.n72 vdd.n71 0.0025
C0 iovdd iovss 0.31051p
C1 vdd iovss 0.24621p
C2 sg13g2_DCNDiode_0.guard iovss 0.27183p $ **FLOATING
.ends

