* NGSPICE file created from OTA_final.ext - technology: ihp-sg13g2

.subckt OTA_final ibias vinn vinp vout vdda vssa
X0 vssa.t16 vssa.t66 vssa.t16 vssa.t4 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X1 w_833_2071.t124 ibias.t12 vssa.t1 vssa.t0 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X2 a_610_6649.t27 vinp.t0 w_833_2071.t22 w_833_2071.t7 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X3 w_833_2071.t40 vinn.t0 vout.t9 w_833_2071.t2 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X4 a_610_6649.t26 vinp.t1 w_833_2071.t17 w_833_2071.t27 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X5 vdda.t68 vdda.t66 vdda.t23 vdda.t0 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X6 vdda.t16 a_610_6649.t28 vout.t0 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X7 w_833_2071.t125 ibias.t13 vssa.t9 vssa.t4 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X8 w_833_2071.t61 w_833_2071.t118 w_833_2071.t61 w_833_2071.t7 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X9 w_833_2071.t25 vinn.t1 vout.t16 w_833_2071.t18 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X10 vdda.t65 vdda.t63 vdda.t1 vdda.t0 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X11 w_833_2071.t10 vinn.t2 vout.t14 w_833_2071.t9 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X12 w_833_2071.t126 vinn.t3 vout.t5 w_833_2071.t16 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X13 w_833_2071.t61 w_833_2071.t116 w_833_2071.t61 w_833_2071.t2 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X14 w_833_2071.t61 w_833_2071.t114 w_833_2071.t61 w_833_2071.t27 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X15 a_610_6649.t24 vinp.t2 w_833_2071.t3 w_833_2071.t43 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X16 vdda.t8 a_610_6649.t9 a_610_6649.t3 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X17 w_833_2071.t55 w_833_2071.t112 w_833_2071.t55 w_833_2071.t18 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X18 vssa.t65 vssa.t63 vssa.t9 vssa.t33 sg13_lv_nmos ad=0.36p pd=2.72u as=0 ps=0 w=1u l=1u
X19 w_833_2071.t55 w_833_2071.t110 w_833_2071.t55 w_833_2071.t16 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X20 ibias.t10 ibias.t11 vssa.t7 vssa.t8 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X21 w_833_2071.t55 w_833_2071.t108 w_833_2071.t55 w_833_2071.t43 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X22 vdda.t18 vdda.t61 vdda.t18 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X23 w_833_2071.t22 vinp.t3 a_610_6649.t20 w_833_2071.t18 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X24 vdda.t5 a_610_6649.t0 a_610_6649.t1 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X25 w_833_2071.t17 vinp.t4 a_610_6649.t27 w_833_2071.t16 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X26 vdda.t23 vdda.t59 vdda.t23 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X27 a_610_6649.t25 vinp.t5 w_833_2071.t53 w_833_2071.t14 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X28 vout.t18 vinn.t4 w_833_2071.t40 w_833_2071.t43 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X29 w_833_2071.t35 vinp.t6 a_610_6649.t19 w_833_2071.t9 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X30 vdda.t13 a_610_6649.t29 vout.t3 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X31 vssa.t16 vssa.t61 vssa.t16 vssa.t6 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X32 vssa.t68 ibias.t14 w_833_2071.t125 vssa.t20 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X33 w_833_2071.t61 w_833_2071.t106 w_833_2071.t61 w_833_2071.t18 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X34 vssa.t21 vssa.t59 vssa.t21 vssa.t8 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X35 vdda.t23 vdda.t57 vdda.t23 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X36 vdda.t7 a_610_6649.t30 vout.t2 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X37 w_833_2071.t61 w_833_2071.t104 w_833_2071.t61 w_833_2071.t16 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X38 vssa.t16 vssa.t57 vssa.t16 vssa.t31 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X39 vssa.t14 ibias.t9 ibias.t10 vssa.t13 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X40 w_833_2071.t61 w_833_2071.t102 w_833_2071.t61 w_833_2071.t43 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X41 vssa.t21 vssa.t55 vssa.t21 vssa.t31 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X42 vdda.t6 a_610_6649.t11 a_610_6649.t7 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X43 vdda.t56 vdda.t54 vdda.t18 vdda.t0 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X44 vssa.t21 vssa.t53 vssa.t21 vssa.t4 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X45 w_833_2071.t122 ibias.t15 vssa.t14 vssa.t0 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X46 vdda.t23 vdda.t52 vdda.t23 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X47 vout.t17 vinn.t5 w_833_2071.t47 w_833_2071.t14 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X48 vdda.t3 a_610_6649.t4 a_610_6649.t5 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X49 w_833_2071.t53 vinp.t7 a_610_6649.t18 w_833_2071.t20 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X50 vssa.t21 vssa.t51 vssa.t21 vssa.t2 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X51 w_833_2071.t123 ibias.t16 vssa.t5 vssa.t4 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X52 vdda.t23 vdda.t50 vdda.t23 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X53 vssa.t45 ibias.t17 w_833_2071.t124 vssa.t11 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X54 vdda.t4 a_610_6649.t31 vout.t1 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X55 vssa.t21 vssa.t49 vssa.t21 vssa.t0 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X56 w_833_2071.t31 vinn.t6 vout.t4 w_833_2071.t9 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X57 vssa.t48 vssa.t46 vssa.t5 vssa.t33 sg13_lv_nmos ad=0.36p pd=2.72u as=0 ps=0 w=1u l=1u
X58 vdda.t18 vdda.t48 vdda.t18 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X59 w_833_2071.t55 w_833_2071.t100 w_833_2071.t55 w_833_2071.t9 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X60 vout.t12 vinn.t7 w_833_2071.t136 w_833_2071.t81 sg13_lv_nmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.5u
X61 vssa.t45 vssa.t44 vssa.t45 vssa.t31 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X62 w_833_2071.t47 vinn.t8 vout.t6 w_833_2071.t20 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X63 vdda.t18 vdda.t46 vdda.t18 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X64 w_833_2071.t1 vinn.t9 vout.t19 w_833_2071.t12 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X65 w_833_2071.t24 vinp.t8 a_610_6649.t26 w_833_2071.t9 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X66 a_610_6649.t23 vinp.t9 w_833_2071.t45 w_833_2071.t5 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X67 vssa.t3 ibias.t18 w_833_2071.t123 vssa.t20 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X68 a_610_6649.t17 vinp.t10 w_833_2071.t21 w_833_2071.t14 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X69 vssa.t16 vssa.t42 vssa.t16 vssa.t20 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X70 w_833_2071.t61 w_833_2071.t98 w_833_2071.t61 w_833_2071.t9 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X71 vssa.t16 vssa.t40 vssa.t16 vssa.t0 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X72 vdda.t18 vdda.t44 vdda.t18 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X73 ibias.t7 ibias.t8 vssa.t68 vssa.t2 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X74 w_833_2071.t55 w_833_2071.t96 w_833_2071.t55 w_833_2071.t14 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X75 a_610_6649.t1 a_610_6649.t8 vdda.t8 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X76 a_610_6649.t14 vinp.t11 w_833_2071.t127 w_833_2071.t81 sg13_lv_nmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.5u
X77 vdda.t18 vdda.t42 vdda.t18 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X78 vssa.t39 vssa.t37 vssa.t16 vssa.t33 sg13_lv_nmos ad=0.36p pd=2.72u as=0 ps=0 w=1u l=1u
X79 vout.t8 vinn.t10 w_833_2071.t15 w_833_2071.t14 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X80 w_833_2071.t13 vinp.t12 a_610_6649.t22 w_833_2071.t12 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X81 vdda.t16 vdda.t40 vdda.t16 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X82 vout.t19 vinn.t11 w_833_2071.t10 w_833_2071.t23 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X83 vout.t15 vinn.t12 w_833_2071.t6 w_833_2071.t5 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X84 a_610_6649.t21 vinp.t13 w_833_2071.t1 w_833_2071.t0 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X85 w_833_2071.t45 vinp.t14 a_610_6649.t25 w_833_2071.t11 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X86 vssa.t12 ibias.t19 w_833_2071.t122 vssa.t11 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X87 w_833_2071.t61 w_833_2071.t94 w_833_2071.t61 w_833_2071.t14 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X88 w_833_2071.t21 vinp.t15 a_610_6649.t24 w_833_2071.t20 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X89 w_833_2071.t42 vinp.t16 a_610_6649.t23 w_833_2071.t33 sg13_lv_nmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.5u
X90 vssa.t10 ibias.t6 ibias.t7 vssa.t6 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X91 vssa.t21 vssa.t35 vssa.t21 vssa.t13 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X92 vdda.t23 vdda.t38 vdda.t23 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X93 a_610_6649.t3 a_610_6649.t2 vdda.t7 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X94 w_833_2071.t55 w_833_2071.t92 w_833_2071.t55 w_833_2071.t20 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X95 vssa.t34 vssa.t32 vssa.t21 vssa.t33 sg13_lv_nmos ad=0.36p pd=2.72u as=0 ps=0 w=1u l=1u
X96 a_610_6649.t5 a_610_6649.t10 vdda.t6 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X97 vdda.t23 vdda.t36 vdda.t23 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X98 vout.t0 a_610_6649.t32 vdda.t5 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X99 w_833_2071.t15 vinn.t13 vout.t18 w_833_2071.t20 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X100 a_610_6649.t22 vinp.t17 w_833_2071.t35 w_833_2071.t23 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X101 vssa.t12 vssa.t30 vssa.t12 vssa.t31 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X102 w_833_2071.t6 vinn.t14 vout.t17 w_833_2071.t11 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X103 vout.t13 vinn.t15 w_833_2071.t13 w_833_2071.t0 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X104 vdda.t13 vdda.t34 vdda.t13 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X105 vout.t11 vinn.t16 w_833_2071.t8 w_833_2071.t7 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X106 vout.t16 vinn.t17 w_833_2071.t129 w_833_2071.t81 sg13_lv_nmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.5u
X107 w_833_2071.t146 vinn.t18 vout.t15 w_833_2071.t33 sg13_lv_nmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.5u
X108 vout.t14 vinn.t19 w_833_2071.t28 w_833_2071.t27 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X109 w_833_2071.t44 vinp.t18 a_610_6649.t21 w_833_2071.t2 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X110 w_833_2071.t61 w_833_2071.t90 w_833_2071.t61 w_833_2071.t20 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X111 w_833_2071.t26 vinn.t20 vout.t10 w_833_2071.t12 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X112 vssa.t16 vssa.t28 vssa.t16 vssa.t8 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X113 vssa.t16 vssa.t26 vssa.t16 vssa.t13 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X114 a_610_6649.t16 vinp.t19 w_833_2071.t48 w_833_2071.t5 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X115 vdda.t23 vdda.t32 vdda.t23 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X116 w_833_2071.t89 w_833_2071.t87 w_833_2071.t55 w_833_2071.t81 sg13_lv_nmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=0.5u
X117 w_833_2071.t55 w_833_2071.t85 w_833_2071.t55 w_833_2071.t12 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X118 ibias.t4 ibias.t5 vssa.t3 vssa.t2 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X119 a_610_6649.t7 a_610_6649.t6 vdda.t4 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X120 vssa.t21 vssa.t24 vssa.t21 vssa.t11 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X121 w_833_2071.t55 w_833_2071.t83 w_833_2071.t55 w_833_2071.t5 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X122 vdda.t23 vdda.t30 vdda.t23 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X123 a_610_6649.t20 vinp.t20 w_833_2071.t140 w_833_2071.t81 sg13_lv_nmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.5u
X124 w_833_2071.t49 vinp.t21 a_610_6649.t15 w_833_2071.t12 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X125 vout.t3 a_610_6649.t33 vdda.t3 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X126 a_610_6649.t13 vinp.t22 w_833_2071.t19 w_833_2071.t7 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X127 a_610_6649.t19 vinp.t23 w_833_2071.t36 w_833_2071.t27 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X128 vssa.t21 vssa.t22 vssa.t21 vssa.t6 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X129 vout.t7 vinn.t21 w_833_2071.t30 w_833_2071.t5 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X130 w_833_2071.t4 vinn.t22 vout.t13 w_833_2071.t2 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X131 w_833_2071.t8 vinn.t23 vout.t12 w_833_2071.t18 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X132 w_833_2071.t28 vinn.t24 vout.t11 w_833_2071.t16 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X133 w_833_2071.t82 w_833_2071.t80 w_833_2071.t61 w_833_2071.t81 sg13_lv_nmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=0.5u
X134 w_833_2071.t61 w_833_2071.t78 w_833_2071.t61 w_833_2071.t12 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X135 vout.t10 vinn.t25 w_833_2071.t31 w_833_2071.t23 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X136 vdda.t18 vdda.t28 vdda.t18 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X137 a_610_6649.t18 vinp.t24 w_833_2071.t44 w_833_2071.t43 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X138 w_833_2071.t48 vinp.t25 a_610_6649.t17 w_833_2071.t11 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X139 a_610_6649.t12 vinp.t26 w_833_2071.t26 w_833_2071.t0 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X140 vout.t2 a_610_6649.t34 vdda.t2 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X141 vssa.t7 ibias.t3 ibias.t4 vssa.t6 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X142 w_833_2071.t61 w_833_2071.t76 w_833_2071.t61 w_833_2071.t5 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X143 w_833_2071.t139 vinp.t27 a_610_6649.t16 w_833_2071.t33 sg13_lv_nmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.5u
X144 vdda.t18 vdda.t26 vdda.t18 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=1u
X145 w_833_2071.t55 w_833_2071.t74 w_833_2071.t55 w_833_2071.t23 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X146 w_833_2071.t55 w_833_2071.t72 w_833_2071.t55 w_833_2071.t0 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X147 w_833_2071.t55 w_833_2071.t70 w_833_2071.t55 w_833_2071.t11 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X148 ibias.t1 ibias.t2 vssa.t10 vssa.t8 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X149 w_833_2071.t55 w_833_2071.t68 w_833_2071.t55 w_833_2071.t33 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X150 vssa.t21 vssa.t19 vssa.t21 vssa.t20 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X151 a_610_6649.t15 vinp.t28 w_833_2071.t24 w_833_2071.t23 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X152 w_833_2071.t19 vinp.t29 a_610_6649.t14 w_833_2071.t18 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X153 vout.t9 vinn.t26 w_833_2071.t49 w_833_2071.t0 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X154 w_833_2071.t36 vinp.t30 a_610_6649.t13 w_833_2071.t16 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X155 w_833_2071.t30 vinn.t27 vout.t8 w_833_2071.t11 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X156 w_833_2071.t34 vinn.t28 vout.t7 w_833_2071.t33 sg13_lv_nmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.5u
X157 vdda.t18 vdda.t24 vdda.t18 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X158 vout.t6 vinn.t29 w_833_2071.t4 w_833_2071.t43 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X159 vdda.t23 vdda.t22 vdda.t23 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X160 vdda.t21 vdda.t19 vdda.t2 vdda.t0 sg13_lv_pmos ad=0.34p pd=2.68u as=0 ps=0 w=1u l=1u
X161 w_833_2071.t61 w_833_2071.t66 w_833_2071.t61 w_833_2071.t23 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X162 vout.t5 vinn.t30 w_833_2071.t25 w_833_2071.t7 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X163 vout.t4 vinn.t31 w_833_2071.t126 w_833_2071.t27 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X164 vssa.t16 vssa.t17 vssa.t16 vssa.t2 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X165 w_833_2071.t61 w_833_2071.t64 w_833_2071.t61 w_833_2071.t11 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X166 w_833_2071.t61 w_833_2071.t62 w_833_2071.t61 w_833_2071.t0 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X167 w_833_2071.t3 vinp.t31 a_610_6649.t12 w_833_2071.t2 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=0.5u
X168 vssa.t1 ibias.t0 ibias.t1 vssa.t13 sg13_lv_nmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X169 w_833_2071.t61 w_833_2071.t60 w_833_2071.t61 w_833_2071.t33 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X170 vout.t1 a_610_6649.t35 vdda.t1 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0.19p ps=1.38u w=1u l=2u
X171 vdda.t18 vdda.t17 vdda.t18 vdda.t0 sg13_lv_pmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X172 vssa.t16 vssa.t15 vssa.t16 vssa.t11 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=2u
X173 w_833_2071.t55 w_833_2071.t58 w_833_2071.t55 w_833_2071.t7 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X174 w_833_2071.t55 w_833_2071.t56 w_833_2071.t55 w_833_2071.t27 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
X175 w_833_2071.t55 w_833_2071.t54 w_833_2071.t55 w_833_2071.t2 sg13_lv_nmos ad=0.19p pd=1.38u as=0 ps=0 w=1u l=0.5u
R0 vssa.t31 vssa.n20 101.591
R1 vssa.t33 vssa.n50 101.591
R2 vssa.t11 vssa.n23 52.335
R3 vssa.n86 vssa.t11 52.335
R4 vssa.n83 vssa.t0 52.335
R5 vssa.t0 vssa.n27 52.335
R6 vssa.t13 vssa.n30 52.335
R7 vssa.n77 vssa.t13 52.335
R8 vssa.n74 vssa.t8 52.335
R9 vssa.t8 vssa.n34 52.335
R10 vssa.t6 vssa.n37 52.335
R11 vssa.n68 vssa.t6 52.335
R12 vssa.n65 vssa.t2 52.335
R13 vssa.t2 vssa.n41 52.335
R14 vssa.t20 vssa.n44 52.335
R15 vssa.n60 vssa.t20 52.335
R16 vssa.n57 vssa.t4 52.335
R17 vssa.t4 vssa.n48 52.335
R18 vssa.n268 vssa.t16 17.1548
R19 vssa.t21 vssa.n166 17.0005
R20 vssa.n251 vssa.n140 17.0005
R21 vssa.n251 vssa.n48 17.0005
R22 vssa.n251 vssa.n60 17.0005
R23 vssa.n251 vssa.n41 17.0005
R24 vssa.n251 vssa.n68 17.0005
R25 vssa.n251 vssa.n34 17.0005
R26 vssa.n251 vssa.n77 17.0005
R27 vssa.n251 vssa.n27 17.0005
R28 vssa.n251 vssa.n86 17.0005
R29 vssa.n251 vssa.n250 17.0005
R30 vssa.n117 vssa.n53 17.0005
R31 vssa.n117 vssa.n50 17.0005
R32 vssa.n117 vssa.n57 17.0005
R33 vssa.n117 vssa.n44 17.0005
R34 vssa.n117 vssa.n65 17.0005
R35 vssa.n117 vssa.n37 17.0005
R36 vssa.n117 vssa.n74 17.0005
R37 vssa.n117 vssa.n30 17.0005
R38 vssa.n117 vssa.n83 17.0005
R39 vssa.n117 vssa.n23 17.0005
R40 vssa.n253 vssa.n117 17.0005
R41 vssa.n117 vssa.n20 17.0005
R42 vssa.n117 vssa.n12 17.0005
R43 vssa.n118 vssa.n117 17.0005
R44 vssa.n140 vssa.n1 17.0005
R45 vssa.n51 vssa.n1 17.0005
R46 vssa.n53 vssa.n1 17.0005
R47 vssa.n50 vssa.n1 17.0005
R48 vssa.n55 vssa.n1 17.0005
R49 vssa.n49 vssa.n1 17.0005
R50 vssa.n56 vssa.n1 17.0005
R51 vssa.n48 vssa.n1 17.0005
R52 vssa.n57 vssa.n1 17.0005
R53 vssa.n47 vssa.n1 17.0005
R54 vssa.n58 vssa.n1 17.0005
R55 vssa.n46 vssa.n1 17.0005
R56 vssa.n59 vssa.n1 17.0005
R57 vssa.n45 vssa.n1 17.0005
R58 vssa.n60 vssa.n1 17.0005
R59 vssa.n44 vssa.n1 17.0005
R60 vssa.n61 vssa.n1 17.0005
R61 vssa.n43 vssa.n1 17.0005
R62 vssa.n63 vssa.n1 17.0005
R63 vssa.n42 vssa.n1 17.0005
R64 vssa.n64 vssa.n1 17.0005
R65 vssa.n41 vssa.n1 17.0005
R66 vssa.n65 vssa.n1 17.0005
R67 vssa.n40 vssa.n1 17.0005
R68 vssa.n66 vssa.n1 17.0005
R69 vssa.n39 vssa.n1 17.0005
R70 vssa.n67 vssa.n1 17.0005
R71 vssa.n38 vssa.n1 17.0005
R72 vssa.n68 vssa.n1 17.0005
R73 vssa.n37 vssa.n1 17.0005
R74 vssa.n69 vssa.n1 17.0005
R75 vssa.n36 vssa.n1 17.0005
R76 vssa.n72 vssa.n1 17.0005
R77 vssa.n35 vssa.n1 17.0005
R78 vssa.n73 vssa.n1 17.0005
R79 vssa.n34 vssa.n1 17.0005
R80 vssa.n74 vssa.n1 17.0005
R81 vssa.n33 vssa.n1 17.0005
R82 vssa.n75 vssa.n1 17.0005
R83 vssa.n32 vssa.n1 17.0005
R84 vssa.n76 vssa.n1 17.0005
R85 vssa.n31 vssa.n1 17.0005
R86 vssa.n77 vssa.n1 17.0005
R87 vssa.n30 vssa.n1 17.0005
R88 vssa.n78 vssa.n1 17.0005
R89 vssa.n29 vssa.n1 17.0005
R90 vssa.n81 vssa.n1 17.0005
R91 vssa.n28 vssa.n1 17.0005
R92 vssa.n82 vssa.n1 17.0005
R93 vssa.n27 vssa.n1 17.0005
R94 vssa.n83 vssa.n1 17.0005
R95 vssa.n26 vssa.n1 17.0005
R96 vssa.n84 vssa.n1 17.0005
R97 vssa.n25 vssa.n1 17.0005
R98 vssa.n85 vssa.n1 17.0005
R99 vssa.n24 vssa.n1 17.0005
R100 vssa.n86 vssa.n1 17.0005
R101 vssa.n23 vssa.n1 17.0005
R102 vssa.n87 vssa.n1 17.0005
R103 vssa.n22 vssa.n1 17.0005
R104 vssa.n90 vssa.n1 17.0005
R105 vssa.n21 vssa.n1 17.0005
R106 vssa.n253 vssa.n1 17.0005
R107 vssa.n20 vssa.n1 17.0005
R108 vssa.n262 vssa.t45 17.0005
R109 vssa.t12 vssa.n162 17.0005
R110 vssa.n254 vssa.n51 17.0005
R111 vssa.n254 vssa.n53 17.0005
R112 vssa.n254 vssa.n50 17.0005
R113 vssa.n254 vssa.n55 17.0005
R114 vssa.n254 vssa.n49 17.0005
R115 vssa.n254 vssa.n56 17.0005
R116 vssa.n254 vssa.n48 17.0005
R117 vssa.n254 vssa.n57 17.0005
R118 vssa.n254 vssa.n47 17.0005
R119 vssa.n254 vssa.n58 17.0005
R120 vssa.n254 vssa.n46 17.0005
R121 vssa.n254 vssa.n59 17.0005
R122 vssa.n254 vssa.n45 17.0005
R123 vssa.n254 vssa.n60 17.0005
R124 vssa.n254 vssa.n44 17.0005
R125 vssa.n254 vssa.n61 17.0005
R126 vssa.n254 vssa.n43 17.0005
R127 vssa.n254 vssa.n63 17.0005
R128 vssa.n254 vssa.n42 17.0005
R129 vssa.n254 vssa.n64 17.0005
R130 vssa.n254 vssa.n41 17.0005
R131 vssa.n254 vssa.n65 17.0005
R132 vssa.n254 vssa.n40 17.0005
R133 vssa.n254 vssa.n66 17.0005
R134 vssa.n254 vssa.n39 17.0005
R135 vssa.n254 vssa.n67 17.0005
R136 vssa.n254 vssa.n38 17.0005
R137 vssa.n254 vssa.n68 17.0005
R138 vssa.n254 vssa.n37 17.0005
R139 vssa.n254 vssa.n69 17.0005
R140 vssa.n254 vssa.n36 17.0005
R141 vssa.n254 vssa.n72 17.0005
R142 vssa.n254 vssa.n35 17.0005
R143 vssa.n254 vssa.n73 17.0005
R144 vssa.n254 vssa.n34 17.0005
R145 vssa.n254 vssa.n74 17.0005
R146 vssa.n254 vssa.n33 17.0005
R147 vssa.n254 vssa.n75 17.0005
R148 vssa.n254 vssa.n32 17.0005
R149 vssa.n254 vssa.n76 17.0005
R150 vssa.n254 vssa.n31 17.0005
R151 vssa.n254 vssa.n77 17.0005
R152 vssa.n254 vssa.n30 17.0005
R153 vssa.n254 vssa.n78 17.0005
R154 vssa.n254 vssa.n29 17.0005
R155 vssa.n254 vssa.n81 17.0005
R156 vssa.n254 vssa.n28 17.0005
R157 vssa.n254 vssa.n82 17.0005
R158 vssa.n254 vssa.n27 17.0005
R159 vssa.n254 vssa.n83 17.0005
R160 vssa.n254 vssa.n26 17.0005
R161 vssa.n254 vssa.n84 17.0005
R162 vssa.n254 vssa.n25 17.0005
R163 vssa.n254 vssa.n85 17.0005
R164 vssa.n254 vssa.n24 17.0005
R165 vssa.n254 vssa.n86 17.0005
R166 vssa.n254 vssa.n23 17.0005
R167 vssa.n254 vssa.n87 17.0005
R168 vssa.n254 vssa.n22 17.0005
R169 vssa.n254 vssa.n90 17.0005
R170 vssa.n254 vssa.n21 17.0005
R171 vssa.n254 vssa.n253 17.0005
R172 vssa.n254 vssa.n20 17.0005
R173 vssa.n254 vssa.n18 17.0005
R174 vssa.n140 vssa.n52 16.9882
R175 vssa.n118 vssa.n52 16.9882
R176 vssa.n116 vssa.n49 13.01
R177 vssa.n116 vssa.n55 13.01
R178 vssa.n119 vssa.n20 12.8328
R179 vssa.n252 vssa.n21 12.8328
R180 vssa.n92 vssa.n21 12.8328
R181 vssa.n121 vssa.n22 12.8328
R182 vssa.n93 vssa.n22 12.8328
R183 vssa.n122 vssa.n23 12.8328
R184 vssa.n94 vssa.n24 12.8328
R185 vssa.n156 vssa.n85 12.8328
R186 vssa.n95 vssa.n25 12.8328
R187 vssa.n155 vssa.n84 12.8328
R188 vssa.n96 vssa.n26 12.8328
R189 vssa.n154 vssa.n83 12.8328
R190 vssa.n97 vssa.n27 12.8328
R191 vssa.n124 vssa.n28 12.8328
R192 vssa.n98 vssa.n28 12.8328
R193 vssa.n125 vssa.n29 12.8328
R194 vssa.n99 vssa.n29 12.8328
R195 vssa.n126 vssa.n30 12.8328
R196 vssa.n100 vssa.n31 12.8328
R197 vssa.n152 vssa.n76 12.8328
R198 vssa.n101 vssa.n32 12.8328
R199 vssa.n151 vssa.n75 12.8328
R200 vssa.n102 vssa.n33 12.8328
R201 vssa.n150 vssa.n74 12.8328
R202 vssa.n103 vssa.n34 12.8328
R203 vssa.n128 vssa.n35 12.8328
R204 vssa.n104 vssa.n35 12.8328
R205 vssa.n129 vssa.n36 12.8328
R206 vssa.n105 vssa.n36 12.8328
R207 vssa.n130 vssa.n37 12.8328
R208 vssa.n106 vssa.n38 12.8328
R209 vssa.n148 vssa.n67 12.8328
R210 vssa.n107 vssa.n39 12.8328
R211 vssa.n147 vssa.n66 12.8328
R212 vssa.n108 vssa.n40 12.8328
R213 vssa.n146 vssa.n65 12.8328
R214 vssa.n109 vssa.n41 12.8328
R215 vssa.n132 vssa.n42 12.8328
R216 vssa.n110 vssa.n42 12.8328
R217 vssa.n133 vssa.n43 12.8328
R218 vssa.n111 vssa.n43 12.8328
R219 vssa.n134 vssa.n44 12.8328
R220 vssa.n112 vssa.n45 12.8328
R221 vssa.n144 vssa.n59 12.8328
R222 vssa.n113 vssa.n46 12.8328
R223 vssa.n143 vssa.n58 12.8328
R224 vssa.n114 vssa.n47 12.8328
R225 vssa.n142 vssa.n57 12.8328
R226 vssa.n115 vssa.n48 12.8328
R227 vssa.n136 vssa.n49 12.8328
R228 vssa.n137 vssa.n50 12.8328
R229 vssa.n138 vssa.n51 12.8328
R230 vssa.n139 vssa.n51 12.8328
R231 vssa.n138 vssa.n53 12.8328
R232 vssa.n137 vssa.n55 12.8328
R233 vssa.n136 vssa.n56 12.8328
R234 vssa.n142 vssa.n47 12.8328
R235 vssa.n143 vssa.n46 12.8328
R236 vssa.n144 vssa.n45 12.8328
R237 vssa.n134 vssa.n61 12.8328
R238 vssa.n133 vssa.n63 12.8328
R239 vssa.n132 vssa.n64 12.8328
R240 vssa.n146 vssa.n40 12.8328
R241 vssa.n147 vssa.n39 12.8328
R242 vssa.n148 vssa.n38 12.8328
R243 vssa.n130 vssa.n69 12.8328
R244 vssa.n129 vssa.n72 12.8328
R245 vssa.n128 vssa.n73 12.8328
R246 vssa.n150 vssa.n33 12.8328
R247 vssa.n151 vssa.n32 12.8328
R248 vssa.n152 vssa.n31 12.8328
R249 vssa.n126 vssa.n78 12.8328
R250 vssa.n125 vssa.n81 12.8328
R251 vssa.n124 vssa.n82 12.8328
R252 vssa.n154 vssa.n26 12.8328
R253 vssa.n155 vssa.n25 12.8328
R254 vssa.n156 vssa.n24 12.8328
R255 vssa.n122 vssa.n87 12.8328
R256 vssa.n121 vssa.n90 12.8328
R257 vssa.n253 vssa.n252 12.8328
R258 vssa.n119 vssa.n118 12.8328
R259 vssa.n140 vssa.n139 12.8328
R260 vssa.n115 vssa.n56 12.8328
R261 vssa.n114 vssa.n58 12.8328
R262 vssa.n113 vssa.n59 12.8328
R263 vssa.n112 vssa.n60 12.8328
R264 vssa.n111 vssa.n61 12.8328
R265 vssa.n110 vssa.n63 12.8328
R266 vssa.n109 vssa.n64 12.8328
R267 vssa.n108 vssa.n66 12.8328
R268 vssa.n107 vssa.n67 12.8328
R269 vssa.n106 vssa.n68 12.8328
R270 vssa.n105 vssa.n69 12.8328
R271 vssa.n104 vssa.n72 12.8328
R272 vssa.n103 vssa.n73 12.8328
R273 vssa.n102 vssa.n75 12.8328
R274 vssa.n101 vssa.n76 12.8328
R275 vssa.n100 vssa.n77 12.8328
R276 vssa.n99 vssa.n78 12.8328
R277 vssa.n98 vssa.n81 12.8328
R278 vssa.n97 vssa.n82 12.8328
R279 vssa.n96 vssa.n84 12.8328
R280 vssa.n95 vssa.n85 12.8328
R281 vssa.n94 vssa.n86 12.8328
R282 vssa.n93 vssa.n87 12.8328
R283 vssa.n92 vssa.n90 12.8328
R284 vssa.n247 vssa.t21 8.49776
R285 vssa.n266 vssa.t16 8.38237
R286 vssa.t45 vssa.n14 8.38237
R287 vssa.n163 vssa.t12 8.38237
R288 vssa.n88 vssa.t14 6.12323
R289 vssa.n79 vssa.t7 6.12323
R290 vssa.n70 vssa.t3 6.12323
R291 vssa.n186 vssa.t1 6.12323
R292 vssa.n188 vssa.t10 6.12323
R293 vssa.n190 vssa.t68 6.12323
R294 vssa.n251 vssa.n120 5.61281
R295 vssa.n117 vssa.n91 5.61281
R296 vssa.n269 vssa.n1 5.61281
R297 vssa.n255 vssa.n254 5.61281
R298 vssa.n220 vssa.t48 5.56245
R299 vssa.n226 vssa.t34 5.56245
R300 vssa.t21 vssa.n171 5.56245
R301 vssa.t21 vssa.n173 5.56245
R302 vssa.t21 vssa.n175 5.56245
R303 vssa.t21 vssa.n177 5.56245
R304 vssa.t21 vssa.n179 5.56245
R305 vssa.t21 vssa.n181 5.56245
R306 vssa.t21 vssa.n183 5.56245
R307 vssa.t21 vssa.n246 5.56245
R308 vssa.t21 vssa.n169 5.56245
R309 vssa.t45 vssa.n261 5.56245
R310 vssa.n184 vssa.t65 5.56245
R311 vssa.n216 vssa.t9 5.56245
R312 vssa.n0 vssa.t39 5.56245
R313 vssa.t16 vssa.n2 5.56245
R314 vssa.t16 vssa.n3 5.56245
R315 vssa.t16 vssa.n4 5.56245
R316 vssa.t16 vssa.n5 5.56245
R317 vssa.t16 vssa.n6 5.56245
R318 vssa.t16 vssa.n7 5.56245
R319 vssa.t16 vssa.n8 5.56245
R320 vssa.t16 vssa.n9 5.56245
R321 vssa.n209 vssa.t16 5.56245
R322 vssa.t12 vssa.n161 5.56245
R323 vssa.n222 vssa.t5 5.56245
R324 vssa.n223 vssa.t46 4.89895
R325 vssa.n167 vssa.t55 4.89895
R326 vssa.n227 vssa.t32 4.89895
R327 vssa.n260 vssa.t44 4.89895
R328 vssa.n217 vssa.t63 4.89895
R329 vssa.n192 vssa.t57 4.89895
R330 vssa.n211 vssa.t37 4.89895
R331 vssa.n160 vssa.t30 4.89895
R332 vssa.n251 vssa.n141 3.30365
R333 vssa.n214 vssa.n117 3.30365
R334 vssa.n287 vssa.n1 3.30365
R335 vssa.n254 vssa.n54 3.30365
R336 vssa.n253 vssa.t31 3.079
R337 vssa.n53 vssa.t33 3.079
R338 vssa.n243 vssa.t24 2.82253
R339 vssa.n241 vssa.t49 2.82253
R340 vssa.n239 vssa.t35 2.82253
R341 vssa.n237 vssa.t59 2.82253
R342 vssa.n235 vssa.t22 2.82253
R343 vssa.n233 vssa.t51 2.82253
R344 vssa.n231 vssa.t19 2.82253
R345 vssa.n229 vssa.t53 2.82253
R346 vssa.n194 vssa.t15 2.82253
R347 vssa.n196 vssa.t40 2.82253
R348 vssa.n198 vssa.t26 2.82253
R349 vssa.n200 vssa.t28 2.82253
R350 vssa.n202 vssa.t61 2.82253
R351 vssa.n204 vssa.t17 2.82253
R352 vssa.n206 vssa.t42 2.82253
R353 vssa.n208 vssa.t66 2.82253
R354 vssa.n251 vssa.n135 2.29333
R355 vssa.n251 vssa.n145 2.29333
R356 vssa.n251 vssa.n131 2.29333
R357 vssa.n251 vssa.n149 2.29333
R358 vssa.n251 vssa.n127 2.29333
R359 vssa.n251 vssa.n153 2.29333
R360 vssa.n251 vssa.n123 2.29333
R361 vssa.n251 vssa.n157 2.29333
R362 vssa.n285 vssa.n1 2.29333
R363 vssa.n283 vssa.n1 2.29333
R364 vssa.n281 vssa.n1 2.29333
R365 vssa.n279 vssa.n1 2.29333
R366 vssa.n277 vssa.n1 2.29333
R367 vssa.n275 vssa.n1 2.29333
R368 vssa.n273 vssa.n1 2.29333
R369 vssa.n271 vssa.n1 2.29333
R370 vssa.n251 vssa.n138 2.0851
R371 vssa.n251 vssa.n137 2.0851
R372 vssa.n251 vssa.n136 2.0851
R373 vssa.n251 vssa.n142 2.0851
R374 vssa.n251 vssa.n143 2.0851
R375 vssa.n251 vssa.n144 2.0851
R376 vssa.n251 vssa.n134 2.0851
R377 vssa.n251 vssa.n133 2.0851
R378 vssa.n251 vssa.n132 2.0851
R379 vssa.n251 vssa.n146 2.0851
R380 vssa.n251 vssa.n147 2.0851
R381 vssa.n251 vssa.n148 2.0851
R382 vssa.n251 vssa.n130 2.0851
R383 vssa.n251 vssa.n129 2.0851
R384 vssa.n251 vssa.n128 2.0851
R385 vssa.n251 vssa.n150 2.0851
R386 vssa.n251 vssa.n151 2.0851
R387 vssa.n251 vssa.n152 2.0851
R388 vssa.n251 vssa.n126 2.0851
R389 vssa.n251 vssa.n125 2.0851
R390 vssa.n251 vssa.n124 2.0851
R391 vssa.n251 vssa.n154 2.0851
R392 vssa.n251 vssa.n155 2.0851
R393 vssa.n251 vssa.n156 2.0851
R394 vssa.n251 vssa.n122 2.0851
R395 vssa.n251 vssa.n121 2.0851
R396 vssa.n252 vssa.n251 2.0851
R397 vssa.n251 vssa.n119 2.0851
R398 vssa.n139 vssa.n117 2.0851
R399 vssa.n117 vssa.n115 2.0851
R400 vssa.n117 vssa.n114 2.0851
R401 vssa.n117 vssa.n113 2.0851
R402 vssa.n117 vssa.n112 2.0851
R403 vssa.n117 vssa.n111 2.0851
R404 vssa.n117 vssa.n110 2.0851
R405 vssa.n117 vssa.n109 2.0851
R406 vssa.n117 vssa.n108 2.0851
R407 vssa.n117 vssa.n107 2.0851
R408 vssa.n117 vssa.n106 2.0851
R409 vssa.n117 vssa.n105 2.0851
R410 vssa.n117 vssa.n104 2.0851
R411 vssa.n117 vssa.n103 2.0851
R412 vssa.n117 vssa.n102 2.0851
R413 vssa.n117 vssa.n101 2.0851
R414 vssa.n117 vssa.n100 2.0851
R415 vssa.n117 vssa.n99 2.0851
R416 vssa.n117 vssa.n98 2.0851
R417 vssa.n117 vssa.n97 2.0851
R418 vssa.n117 vssa.n96 2.0851
R419 vssa.n117 vssa.n95 2.0851
R420 vssa.n117 vssa.n94 2.0851
R421 vssa.n117 vssa.n93 2.0851
R422 vssa.n117 vssa.n92 2.0851
R423 vssa.n117 vssa.n116 1.9965
R424 vssa vssa.n288 1.46167
R425 vssa.n249 vssa.n248 1.073
R426 vssa.n259 vssa.n13 1.073
R427 vssa.n267 vssa.n10 1.073
R428 vssa.n159 vssa.n17 1.073
R429 vssa.n13 vssa.n11 1.06612
R430 vssa.n256 vssa.n17 1.06612
R431 vssa.n261 vssa.n260 0.975229
R432 vssa.n161 vssa.n160 0.975229
R433 vssa.n223 vssa.n222 0.974882
R434 vssa.n227 vssa.n226 0.974882
R435 vssa.n217 vssa.n216 0.974882
R436 vssa.n191 vssa.n117 0.96926
R437 vssa.n189 vssa.n117 0.96926
R438 vssa.n187 vssa.n117 0.96926
R439 vssa.n185 vssa.n117 0.96926
R440 vssa.n254 vssa.n62 0.96926
R441 vssa.n254 vssa.n71 0.96926
R442 vssa.n254 vssa.n80 0.96926
R443 vssa.n254 vssa.n89 0.96926
R444 vssa.n247 vssa.n167 0.856338
R445 vssa.n186 vssa.n185 0.853661
R446 vssa.n188 vssa.n187 0.853661
R447 vssa.n190 vssa.n189 0.853661
R448 vssa.n215 vssa.n191 0.853661
R449 vssa.n89 vssa.n88 0.853661
R450 vssa.n80 vssa.n79 0.853661
R451 vssa.n71 vssa.n70 0.853661
R452 vssa.n221 vssa.n62 0.853661
R453 vssa.n164 vssa.n163 0.841843
R454 vssa.n266 vssa.n265 0.841555
R455 vssa.n258 vssa.n14 0.841555
R456 vssa.n243 vssa.n242 0.803704
R457 vssa.n241 vssa.n240 0.803704
R458 vssa.n239 vssa.n238 0.803704
R459 vssa.n237 vssa.n236 0.803704
R460 vssa.n235 vssa.n234 0.803704
R461 vssa.n233 vssa.n232 0.803704
R462 vssa.n231 vssa.n230 0.803704
R463 vssa.n229 vssa.n228 0.803704
R464 vssa.n195 vssa.n194 0.803704
R465 vssa.n197 vssa.n196 0.803704
R466 vssa.n199 vssa.n198 0.803704
R467 vssa.n201 vssa.n200 0.803704
R468 vssa.n203 vssa.n202 0.803704
R469 vssa.n205 vssa.n204 0.803704
R470 vssa.n207 vssa.n206 0.803704
R471 vssa.n210 vssa.n208 0.803704
R472 vssa.n244 vssa.n243 0.802423
R473 vssa.n242 vssa.n241 0.802423
R474 vssa.n240 vssa.n239 0.802423
R475 vssa.n238 vssa.n237 0.802423
R476 vssa.n236 vssa.n235 0.802423
R477 vssa.n234 vssa.n233 0.802423
R478 vssa.n232 vssa.n231 0.802423
R479 vssa.n230 vssa.n229 0.802423
R480 vssa.n194 vssa.n193 0.802423
R481 vssa.n196 vssa.n195 0.802423
R482 vssa.n198 vssa.n197 0.802423
R483 vssa.n200 vssa.n199 0.802423
R484 vssa.n202 vssa.n201 0.802423
R485 vssa.n204 vssa.n203 0.802423
R486 vssa.n206 vssa.n205 0.802423
R487 vssa.n208 vssa.n207 0.802423
R488 vssa.n166 vssa.n158 0.763625
R489 vssa.n263 vssa.n262 0.75675
R490 vssa.n162 vssa.n16 0.75675
R491 vssa.n185 vssa.n15 0.72267
R492 vssa.n187 vssa.n186 0.72267
R493 vssa.n189 vssa.n188 0.72267
R494 vssa.n191 vssa.n190 0.72267
R495 vssa.n89 vssa.n19 0.72267
R496 vssa.n88 vssa.n80 0.72267
R497 vssa.n79 vssa.n71 0.72267
R498 vssa.n70 vssa.n62 0.72267
R499 vssa.n269 vssa.n268 0.633808
R500 vssa.n226 vssa.n225 0.565495
R501 vssa.n171 vssa.n170 0.565149
R502 vssa.n173 vssa.n172 0.565149
R503 vssa.n175 vssa.n174 0.565149
R504 vssa.n177 vssa.n176 0.565149
R505 vssa.n179 vssa.n178 0.565149
R506 vssa.n181 vssa.n180 0.565149
R507 vssa.n183 vssa.n182 0.565149
R508 vssa.n246 vssa.n245 0.565149
R509 vssa.n220 vssa.n219 0.562058
R510 vssa.n261 vssa.n15 0.562058
R511 vssa.n213 vssa.n184 0.562058
R512 vssa.n288 vssa.n0 0.562058
R513 vssa.n270 vssa.n9 0.562058
R514 vssa.n161 vssa.n19 0.562058
R515 vssa.n284 vssa.n2 0.561712
R516 vssa.n282 vssa.n3 0.561712
R517 vssa.n280 vssa.n4 0.561712
R518 vssa.n278 vssa.n5 0.561712
R519 vssa.n276 vssa.n6 0.561712
R520 vssa.n274 vssa.n7 0.561712
R521 vssa.n272 vssa.n8 0.561712
R522 vssa.n230 vssa.n171 0.50362
R523 vssa.n232 vssa.n173 0.50362
R524 vssa.n234 vssa.n175 0.50362
R525 vssa.n236 vssa.n177 0.50362
R526 vssa.n238 vssa.n179 0.50362
R527 vssa.n240 vssa.n181 0.50362
R528 vssa.n242 vssa.n183 0.50362
R529 vssa.n246 vssa.n244 0.50362
R530 vssa.n228 vssa.n169 0.50362
R531 vssa.n207 vssa.n2 0.50362
R532 vssa.n205 vssa.n3 0.50362
R533 vssa.n203 vssa.n4 0.50362
R534 vssa.n201 vssa.n5 0.50362
R535 vssa.n199 vssa.n6 0.50362
R536 vssa.n197 vssa.n7 0.50362
R537 vssa.n195 vssa.n8 0.50362
R538 vssa.n210 vssa.n209 0.50362
R539 vssa.n224 vssa.n220 0.503274
R540 vssa.n218 vssa.n184 0.503274
R541 vssa.n212 vssa.n0 0.503274
R542 vssa.n193 vssa.n9 0.503274
R543 vssa.n216 vssa 0.500183
R544 vssa.n169 vssa 0.499837
R545 vssa.n182 vssa.n157 0.49086
R546 vssa.n180 vssa.n123 0.49086
R547 vssa.n178 vssa.n153 0.49086
R548 vssa.n176 vssa.n127 0.49086
R549 vssa.n174 vssa.n149 0.49086
R550 vssa.n172 vssa.n131 0.49086
R551 vssa.n170 vssa.n145 0.49086
R552 vssa.n168 vssa.n135 0.49086
R553 vssa.n272 vssa.n271 0.49086
R554 vssa.n274 vssa.n273 0.49086
R555 vssa.n276 vssa.n275 0.49086
R556 vssa.n278 vssa.n277 0.49086
R557 vssa.n280 vssa.n279 0.49086
R558 vssa.n282 vssa.n281 0.49086
R559 vssa.n284 vssa.n283 0.49086
R560 vssa.n286 vssa.n285 0.49086
R561 vssa.n224 vssa.n223 0.472454
R562 vssa.n244 vssa.n167 0.472454
R563 vssa.n228 vssa.n227 0.472454
R564 vssa.n218 vssa.n217 0.472454
R565 vssa.n193 vssa.n192 0.472454
R566 vssa.n212 vssa.n211 0.472454
R567 vssa.n209 vssa 0.472337
R568 vssa.n211 vssa.n210 0.472107
R569 vssa.n260 vssa.n259 0.444607
R570 vssa.n192 vssa.n10 0.444607
R571 vssa.n160 vssa.n159 0.444607
R572 vssa.n222 vssa 0.431433
R573 vssa.n248 vssa.n166 0.419875
R574 vssa.n262 vssa.n13 0.419875
R575 vssa.n162 vssa.n17 0.419875
R576 vssa.n245 vssa.n157 0.363944
R577 vssa.n182 vssa.n123 0.363944
R578 vssa.n180 vssa.n153 0.363944
R579 vssa.n178 vssa.n127 0.363944
R580 vssa.n176 vssa.n149 0.363944
R581 vssa.n174 vssa.n131 0.363944
R582 vssa.n172 vssa.n145 0.363944
R583 vssa.n170 vssa.n135 0.363944
R584 vssa.n271 vssa.n270 0.363944
R585 vssa.n273 vssa.n272 0.363944
R586 vssa.n275 vssa.n274 0.363944
R587 vssa.n277 vssa.n276 0.363944
R588 vssa.n279 vssa.n278 0.363944
R589 vssa.n281 vssa.n280 0.363944
R590 vssa.n283 vssa.n282 0.363944
R591 vssa.n285 vssa.n284 0.363944
R592 vssa.n267 vssa.n266 0.300142
R593 vssa.n14 vssa.n13 0.300142
R594 vssa.n163 vssa.n17 0.300142
R595 vssa.n264 vssa.n263 0.282375
R596 vssa.n257 vssa.n16 0.282375
R597 vssa.n168 vssa.n141 0.254033
R598 vssa.n215 vssa.n214 0.254033
R599 vssa.n287 vssa.n286 0.254033
R600 vssa.n221 vssa.n54 0.254033
R601 vssa.n245 vssa.n120 0.250092
R602 vssa.n91 vssa.n15 0.250092
R603 vssa.n270 vssa.n269 0.250092
R604 vssa.n255 vssa.n19 0.250092
R605 vssa.n225 vssa.n141 0.247939
R606 vssa.n214 vssa.n213 0.247939
R607 vssa.n288 vssa.n287 0.247939
R608 vssa.n219 vssa.n54 0.247939
R609 vssa.n249 vssa.n120 0.242419
R610 vssa.n91 vssa.n11 0.242419
R611 vssa.n256 vssa.n255 0.242419
R612 vssa.n165 vssa.n158 0.23425
R613 vssa.n268 vssa.n267 0.19155
R614 vssa.n264 vssa.n11 0.172375
R615 vssa.n219 vssa.n218 0.172375
R616 vssa.n213 vssa.n212 0.172375
R617 vssa.n257 vssa.n256 0.172375
R618 vssa.n248 vssa.n247 0.145405
R619 vssa vssa.n221 0.131125
R620 vssa.n225 vssa.n224 0.12425
R621 vssa.n249 vssa.n165 0.12425
R622 vssa.n265 vssa.n264 0.0931675
R623 vssa.n258 vssa.n257 0.0931675
R624 vssa.n165 vssa.n164 0.0686545
R625 vssa vssa.n168 0.0658125
R626 vssa vssa.n215 0.062375
R627 vssa.n286 vssa 0.062375
R628 vssa.n259 vssa.n258 0.0119941
R629 vssa.n265 vssa.n10 0.0119941
R630 vssa.n164 vssa.n159 0.0111992
R631 vssa.n250 vssa.n158 0.00783333
R632 vssa.n250 vssa.n249 0.00783333
R633 vssa.n263 vssa.n12 0.00783333
R634 vssa.n12 vssa.n11 0.00783333
R635 vssa.n18 vssa.n16 0.00783333
R636 vssa.n256 vssa.n18 0.00783333
R637 vssa.n254 vssa.n52 0.00738195
R638 ibias.n22 ibias.n0 10.8172
R639 ibias.n22 ibias.n21 9.37277
R640 ibias.n15 ibias.t10 5.6534
R641 ibias.n20 ibias.t4 5.6534
R642 ibias.n10 ibias.t7 5.6534
R643 ibias.n5 ibias.t1 5.6534
R644 ibias.n11 ibias.t16 4.42794
R645 ibias.n13 ibias.t19 4.42666
R646 ibias.n3 ibias.t17 4.42666
R647 ibias.n1 ibias.t13 4.42557
R648 ibias ibias.n22 3.81636
R649 ibias.n21 ibias.n10 3.73245
R650 ibias.n5 ibias.n0 3.73245
R651 ibias.n15 ibias.n0 3.04514
R652 ibias.n21 ibias.n20 3.04514
R653 ibias.n2 ibias.t8 2.82253
R654 ibias.n1 ibias.t14 2.82253
R655 ibias.n13 ibias.t15 2.82253
R656 ibias.n14 ibias.t9 2.82253
R657 ibias.n12 ibias.t5 2.82253
R658 ibias.n11 ibias.t18 2.82253
R659 ibias.n17 ibias.t11 2.82253
R660 ibias.n18 ibias.t3 2.82253
R661 ibias.n7 ibias.t2 2.82253
R662 ibias.n8 ibias.t6 2.82253
R663 ibias.n3 ibias.t12 2.82253
R664 ibias.n4 ibias.t0 2.82253
R665 ibias.n2 ibias.n1 1.60563
R666 ibias.n14 ibias.n13 1.60563
R667 ibias.n12 ibias.n11 1.60563
R668 ibias.n18 ibias.n17 1.60563
R669 ibias.n8 ibias.n7 1.60563
R670 ibias.n4 ibias.n3 1.60563
R671 ibias.n16 ibias.n14 0.704016
R672 ibias.n19 ibias.n18 0.704016
R673 ibias.n9 ibias.n8 0.704016
R674 ibias.n6 ibias.n4 0.704016
R675 ibias.n9 ibias.n2 0.702736
R676 ibias.n19 ibias.n12 0.702736
R677 ibias.n17 ibias.n16 0.702736
R678 ibias.n7 ibias.n6 0.702736
R679 ibias.n16 ibias.n15 0.26531
R680 ibias.n20 ibias.n19 0.26531
R681 ibias.n10 ibias.n9 0.26531
R682 ibias.n6 ibias.n5 0.26531
R683 w_833_2071.n296 w_833_2071.n34 60.1886
R684 w_833_2071.n279 w_833_2071.t33 56.4268
R685 w_833_2071.n280 w_833_2071.n53 56.4268
R686 w_833_2071.n281 w_833_2071.n52 56.4268
R687 w_833_2071.n277 w_833_2071.n6 56.4268
R688 w_833_2071.n276 w_833_2071.n8 56.4268
R689 w_833_2071.n275 w_833_2071.n9 56.4268
R690 w_833_2071.n284 w_833_2071.n49 56.4268
R691 w_833_2071.n285 w_833_2071.n48 56.4268
R692 w_833_2071.n273 w_833_2071.n14 56.4268
R693 w_833_2071.n286 w_833_2071.n47 56.4268
R694 w_833_2071.n272 w_833_2071.n15 56.4268
R695 w_833_2071.n271 w_833_2071.n16 56.4268
R696 w_833_2071.n288 w_833_2071.n45 56.4268
R697 w_833_2071.n289 w_833_2071.n44 56.4268
R698 w_833_2071.n290 w_833_2071.n43 56.4268
R699 w_833_2071.n267 w_833_2071.n19 56.4268
R700 w_833_2071.n266 w_833_2071.n20 56.4268
R701 w_833_2071.t9 w_833_2071.n41 56.4268
R702 w_833_2071.n265 w_833_2071.n21 56.4268
R703 w_833_2071.n292 w_833_2071.n38 56.4268
R704 w_833_2071.n293 w_833_2071.n37 56.4268
R705 w_833_2071.n263 w_833_2071.n23 56.4268
R706 w_833_2071.n262 w_833_2071.n25 56.4268
R707 w_833_2071.n261 w_833_2071.n26 56.4268
R708 w_833_2071.n297 w_833_2071.n31 56.4268
R709 w_833_2071.n298 w_833_2071.n30 56.4268
R710 w_833_2071.n294 w_833_2071.t16 52.6651
R711 w_833_2071.t14 w_833_2071.n50 48.9033
R712 w_833_2071.n269 w_833_2071.t0 48.9033
R713 w_833_2071.t81 w_833_2071.n28 48.9033
R714 w_833_2071.n282 w_833_2071.t11 45.1416
R715 w_833_2071.t12 w_833_2071.n18 45.1416
R716 w_833_2071.n260 w_833_2071.t18 45.1416
R717 w_833_2071.t7 w_833_2071.n35 41.3798
R718 w_833_2071.t5 w_833_2071.n5 37.6181
R719 w_833_2071.n291 w_833_2071.t23 37.6181
R720 w_833_2071.n274 w_833_2071.t20 33.8563
R721 w_833_2071.t2 w_833_2071.n46 33.8563
R722 w_833_2071.t27 w_833_2071.n22 30.0945
R723 w_833_2071.n264 w_833_2071.t27 26.3328
R724 w_833_2071.t20 w_833_2071.n10 22.571
R725 w_833_2071.n287 w_833_2071.t2 22.571
R726 w_833_2071.n278 w_833_2071.t5 18.8093
R727 w_833_2071.t23 w_833_2071.n42 18.8093
R728 w_833_2071.n56 w_833_2071.t33 17.3178
R729 w_833_2071.t55 w_833_2071.n218 17.0005
R730 w_833_2071.n186 w_833_2071.t61 17.0005
R731 w_833_2071.n89 w_833_2071.n30 17.0005
R732 w_833_2071.n89 w_833_2071.n28 17.0005
R733 w_833_2071.n89 w_833_2071.n31 17.0005
R734 w_833_2071.n89 w_833_2071.n27 17.0005
R735 w_833_2071.n89 w_833_2071.n34 17.0005
R736 w_833_2071.n89 w_833_2071.n26 17.0005
R737 w_833_2071.n89 w_833_2071.n35 17.0005
R738 w_833_2071.n89 w_833_2071.n25 17.0005
R739 w_833_2071.n89 w_833_2071.n36 17.0005
R740 w_833_2071.n89 w_833_2071.n23 17.0005
R741 w_833_2071.n89 w_833_2071.n37 17.0005
R742 w_833_2071.n89 w_833_2071.n22 17.0005
R743 w_833_2071.n89 w_833_2071.n38 17.0005
R744 w_833_2071.n89 w_833_2071.n21 17.0005
R745 w_833_2071.n89 w_833_2071.n41 17.0005
R746 w_833_2071.n89 w_833_2071.n20 17.0005
R747 w_833_2071.n89 w_833_2071.n42 17.0005
R748 w_833_2071.n89 w_833_2071.n19 17.0005
R749 w_833_2071.n134 w_833_2071.n89 17.0005
R750 w_833_2071.n89 w_833_2071.n29 17.0005
R751 w_833_2071.n322 w_833_2071.n89 17.0005
R752 w_833_2071.n89 w_833_2071.t33 17.0005
R753 w_833_2071.n89 w_833_2071.n53 17.0005
R754 w_833_2071.n89 w_833_2071.n5 17.0005
R755 w_833_2071.n89 w_833_2071.n52 17.0005
R756 w_833_2071.n89 w_833_2071.n6 17.0005
R757 w_833_2071.n89 w_833_2071.n51 17.0005
R758 w_833_2071.n89 w_833_2071.n8 17.0005
R759 w_833_2071.n89 w_833_2071.n50 17.0005
R760 w_833_2071.n89 w_833_2071.n9 17.0005
R761 w_833_2071.n89 w_833_2071.n49 17.0005
R762 w_833_2071.n89 w_833_2071.n10 17.0005
R763 w_833_2071.n89 w_833_2071.n48 17.0005
R764 w_833_2071.n89 w_833_2071.n14 17.0005
R765 w_833_2071.n89 w_833_2071.n47 17.0005
R766 w_833_2071.n89 w_833_2071.n15 17.0005
R767 w_833_2071.n89 w_833_2071.n46 17.0005
R768 w_833_2071.n89 w_833_2071.n16 17.0005
R769 w_833_2071.n89 w_833_2071.n45 17.0005
R770 w_833_2071.n89 w_833_2071.n17 17.0005
R771 w_833_2071.n89 w_833_2071.n44 17.0005
R772 w_833_2071.n89 w_833_2071.n18 17.0005
R773 w_833_2071.n89 w_833_2071.n43 17.0005
R774 w_833_2071.n196 w_833_2071.n29 17.0005
R775 w_833_2071.n196 w_833_2071.n30 17.0005
R776 w_833_2071.n196 w_833_2071.n28 17.0005
R777 w_833_2071.n196 w_833_2071.n31 17.0005
R778 w_833_2071.n196 w_833_2071.n27 17.0005
R779 w_833_2071.n196 w_833_2071.n34 17.0005
R780 w_833_2071.n196 w_833_2071.n26 17.0005
R781 w_833_2071.n196 w_833_2071.n35 17.0005
R782 w_833_2071.n196 w_833_2071.n25 17.0005
R783 w_833_2071.n196 w_833_2071.n36 17.0005
R784 w_833_2071.n196 w_833_2071.n23 17.0005
R785 w_833_2071.n196 w_833_2071.n37 17.0005
R786 w_833_2071.n196 w_833_2071.n22 17.0005
R787 w_833_2071.n196 w_833_2071.n38 17.0005
R788 w_833_2071.n196 w_833_2071.n21 17.0005
R789 w_833_2071.n196 w_833_2071.n41 17.0005
R790 w_833_2071.n196 w_833_2071.n20 17.0005
R791 w_833_2071.n196 w_833_2071.n42 17.0005
R792 w_833_2071.n196 w_833_2071.n19 17.0005
R793 w_833_2071.n196 w_833_2071.n43 17.0005
R794 w_833_2071.n196 w_833_2071.n18 17.0005
R795 w_833_2071.n196 w_833_2071.n44 17.0005
R796 w_833_2071.n196 w_833_2071.n17 17.0005
R797 w_833_2071.n196 w_833_2071.n45 17.0005
R798 w_833_2071.n196 w_833_2071.n16 17.0005
R799 w_833_2071.n196 w_833_2071.n46 17.0005
R800 w_833_2071.n196 w_833_2071.n15 17.0005
R801 w_833_2071.n196 w_833_2071.n47 17.0005
R802 w_833_2071.n196 w_833_2071.n14 17.0005
R803 w_833_2071.n196 w_833_2071.n48 17.0005
R804 w_833_2071.n196 w_833_2071.n10 17.0005
R805 w_833_2071.n196 w_833_2071.n49 17.0005
R806 w_833_2071.n196 w_833_2071.n9 17.0005
R807 w_833_2071.n196 w_833_2071.n50 17.0005
R808 w_833_2071.n196 w_833_2071.n8 17.0005
R809 w_833_2071.n196 w_833_2071.n51 17.0005
R810 w_833_2071.n196 w_833_2071.n6 17.0005
R811 w_833_2071.n196 w_833_2071.n52 17.0005
R812 w_833_2071.n196 w_833_2071.n5 17.0005
R813 w_833_2071.n196 w_833_2071.n53 17.0005
R814 w_833_2071.n196 w_833_2071.t33 17.0005
R815 w_833_2071.n322 w_833_2071.n196 17.0005
R816 w_833_2071.n88 w_833_2071.n29 17.0005
R817 w_833_2071.n88 w_833_2071.n30 17.0005
R818 w_833_2071.n88 w_833_2071.n28 17.0005
R819 w_833_2071.n88 w_833_2071.n31 17.0005
R820 w_833_2071.n88 w_833_2071.n27 17.0005
R821 w_833_2071.n88 w_833_2071.n34 17.0005
R822 w_833_2071.n88 w_833_2071.n26 17.0005
R823 w_833_2071.n88 w_833_2071.n35 17.0005
R824 w_833_2071.n88 w_833_2071.n25 17.0005
R825 w_833_2071.n88 w_833_2071.n36 17.0005
R826 w_833_2071.n88 w_833_2071.n23 17.0005
R827 w_833_2071.n88 w_833_2071.n37 17.0005
R828 w_833_2071.n88 w_833_2071.n22 17.0005
R829 w_833_2071.n88 w_833_2071.n38 17.0005
R830 w_833_2071.n88 w_833_2071.n21 17.0005
R831 w_833_2071.n88 w_833_2071.n41 17.0005
R832 w_833_2071.n88 w_833_2071.n20 17.0005
R833 w_833_2071.n88 w_833_2071.n42 17.0005
R834 w_833_2071.n88 w_833_2071.n19 17.0005
R835 w_833_2071.n88 w_833_2071.n43 17.0005
R836 w_833_2071.n88 w_833_2071.n18 17.0005
R837 w_833_2071.n88 w_833_2071.n44 17.0005
R838 w_833_2071.n88 w_833_2071.n17 17.0005
R839 w_833_2071.n88 w_833_2071.n45 17.0005
R840 w_833_2071.n88 w_833_2071.n16 17.0005
R841 w_833_2071.n88 w_833_2071.n46 17.0005
R842 w_833_2071.n88 w_833_2071.n15 17.0005
R843 w_833_2071.n88 w_833_2071.n47 17.0005
R844 w_833_2071.n88 w_833_2071.n14 17.0005
R845 w_833_2071.n88 w_833_2071.n48 17.0005
R846 w_833_2071.n88 w_833_2071.n10 17.0005
R847 w_833_2071.n88 w_833_2071.n49 17.0005
R848 w_833_2071.n88 w_833_2071.n9 17.0005
R849 w_833_2071.n88 w_833_2071.n50 17.0005
R850 w_833_2071.n88 w_833_2071.n8 17.0005
R851 w_833_2071.n88 w_833_2071.n51 17.0005
R852 w_833_2071.n88 w_833_2071.n6 17.0005
R853 w_833_2071.n88 w_833_2071.n52 17.0005
R854 w_833_2071.n88 w_833_2071.n5 17.0005
R855 w_833_2071.n88 w_833_2071.n53 17.0005
R856 w_833_2071.n88 w_833_2071.t33 17.0005
R857 w_833_2071.n322 w_833_2071.n88 17.0005
R858 w_833_2071.n323 w_833_2071.n29 17.0005
R859 w_833_2071.n323 w_833_2071.n30 17.0005
R860 w_833_2071.n323 w_833_2071.n28 17.0005
R861 w_833_2071.n323 w_833_2071.n31 17.0005
R862 w_833_2071.n323 w_833_2071.n27 17.0005
R863 w_833_2071.n323 w_833_2071.n34 17.0005
R864 w_833_2071.n323 w_833_2071.n26 17.0005
R865 w_833_2071.n323 w_833_2071.n35 17.0005
R866 w_833_2071.n323 w_833_2071.n25 17.0005
R867 w_833_2071.n323 w_833_2071.n36 17.0005
R868 w_833_2071.n323 w_833_2071.n23 17.0005
R869 w_833_2071.n323 w_833_2071.n37 17.0005
R870 w_833_2071.n323 w_833_2071.n22 17.0005
R871 w_833_2071.n323 w_833_2071.n38 17.0005
R872 w_833_2071.n323 w_833_2071.n21 17.0005
R873 w_833_2071.n323 w_833_2071.n41 17.0005
R874 w_833_2071.n323 w_833_2071.n20 17.0005
R875 w_833_2071.n323 w_833_2071.n42 17.0005
R876 w_833_2071.n323 w_833_2071.n19 17.0005
R877 w_833_2071.n323 w_833_2071.n43 17.0005
R878 w_833_2071.n323 w_833_2071.n18 17.0005
R879 w_833_2071.n323 w_833_2071.n44 17.0005
R880 w_833_2071.n323 w_833_2071.n17 17.0005
R881 w_833_2071.n323 w_833_2071.n45 17.0005
R882 w_833_2071.n323 w_833_2071.n16 17.0005
R883 w_833_2071.n323 w_833_2071.n46 17.0005
R884 w_833_2071.n323 w_833_2071.n15 17.0005
R885 w_833_2071.n323 w_833_2071.n47 17.0005
R886 w_833_2071.n323 w_833_2071.n14 17.0005
R887 w_833_2071.n323 w_833_2071.n48 17.0005
R888 w_833_2071.n323 w_833_2071.n10 17.0005
R889 w_833_2071.n323 w_833_2071.n49 17.0005
R890 w_833_2071.n323 w_833_2071.n9 17.0005
R891 w_833_2071.n323 w_833_2071.n50 17.0005
R892 w_833_2071.n323 w_833_2071.n8 17.0005
R893 w_833_2071.n323 w_833_2071.n51 17.0005
R894 w_833_2071.n323 w_833_2071.n6 17.0005
R895 w_833_2071.n323 w_833_2071.n52 17.0005
R896 w_833_2071.n323 w_833_2071.n5 17.0005
R897 w_833_2071.n323 w_833_2071.n53 17.0005
R898 w_833_2071.n323 w_833_2071.t33 17.0005
R899 w_833_2071.n323 w_833_2071.n322 17.0005
R900 w_833_2071.n321 w_833_2071.n29 17.0005
R901 w_833_2071.n321 w_833_2071.n30 17.0005
R902 w_833_2071.n321 w_833_2071.n28 17.0005
R903 w_833_2071.n321 w_833_2071.n31 17.0005
R904 w_833_2071.n321 w_833_2071.n27 17.0005
R905 w_833_2071.n321 w_833_2071.n34 17.0005
R906 w_833_2071.n321 w_833_2071.n26 17.0005
R907 w_833_2071.n321 w_833_2071.n35 17.0005
R908 w_833_2071.n321 w_833_2071.n25 17.0005
R909 w_833_2071.n321 w_833_2071.n36 17.0005
R910 w_833_2071.n321 w_833_2071.n23 17.0005
R911 w_833_2071.n321 w_833_2071.n37 17.0005
R912 w_833_2071.n321 w_833_2071.n22 17.0005
R913 w_833_2071.n321 w_833_2071.n38 17.0005
R914 w_833_2071.n321 w_833_2071.n21 17.0005
R915 w_833_2071.n321 w_833_2071.n41 17.0005
R916 w_833_2071.n321 w_833_2071.n20 17.0005
R917 w_833_2071.n321 w_833_2071.n42 17.0005
R918 w_833_2071.n321 w_833_2071.n19 17.0005
R919 w_833_2071.n321 w_833_2071.n43 17.0005
R920 w_833_2071.n321 w_833_2071.n18 17.0005
R921 w_833_2071.n321 w_833_2071.n44 17.0005
R922 w_833_2071.n321 w_833_2071.n17 17.0005
R923 w_833_2071.n321 w_833_2071.n45 17.0005
R924 w_833_2071.n321 w_833_2071.n16 17.0005
R925 w_833_2071.n321 w_833_2071.n46 17.0005
R926 w_833_2071.n321 w_833_2071.n15 17.0005
R927 w_833_2071.n321 w_833_2071.n47 17.0005
R928 w_833_2071.n321 w_833_2071.n14 17.0005
R929 w_833_2071.n321 w_833_2071.n48 17.0005
R930 w_833_2071.n321 w_833_2071.n10 17.0005
R931 w_833_2071.n321 w_833_2071.n49 17.0005
R932 w_833_2071.n321 w_833_2071.n9 17.0005
R933 w_833_2071.n321 w_833_2071.n50 17.0005
R934 w_833_2071.n321 w_833_2071.n8 17.0005
R935 w_833_2071.n321 w_833_2071.n51 17.0005
R936 w_833_2071.n321 w_833_2071.n6 17.0005
R937 w_833_2071.n321 w_833_2071.n52 17.0005
R938 w_833_2071.n321 w_833_2071.n5 17.0005
R939 w_833_2071.n321 w_833_2071.n53 17.0005
R940 w_833_2071.n321 w_833_2071.t33 17.0005
R941 w_833_2071.n322 w_833_2071.n321 17.0005
R942 w_833_2071.n299 w_833_2071.n279 17.0005
R943 w_833_2071.n299 w_833_2071.n280 17.0005
R944 w_833_2071.n299 w_833_2071.n278 17.0005
R945 w_833_2071.n299 w_833_2071.n281 17.0005
R946 w_833_2071.n299 w_833_2071.n277 17.0005
R947 w_833_2071.n299 w_833_2071.n282 17.0005
R948 w_833_2071.n299 w_833_2071.n276 17.0005
R949 w_833_2071.n299 w_833_2071.n283 17.0005
R950 w_833_2071.n299 w_833_2071.n275 17.0005
R951 w_833_2071.n299 w_833_2071.n284 17.0005
R952 w_833_2071.n299 w_833_2071.n274 17.0005
R953 w_833_2071.n299 w_833_2071.n285 17.0005
R954 w_833_2071.n299 w_833_2071.n273 17.0005
R955 w_833_2071.n299 w_833_2071.n286 17.0005
R956 w_833_2071.n299 w_833_2071.n272 17.0005
R957 w_833_2071.n299 w_833_2071.n287 17.0005
R958 w_833_2071.n299 w_833_2071.n271 17.0005
R959 w_833_2071.n299 w_833_2071.n288 17.0005
R960 w_833_2071.n299 w_833_2071.n269 17.0005
R961 w_833_2071.n299 w_833_2071.n289 17.0005
R962 w_833_2071.n299 w_833_2071.n268 17.0005
R963 w_833_2071.n299 w_833_2071.n290 17.0005
R964 w_833_2071.n299 w_833_2071.n267 17.0005
R965 w_833_2071.n299 w_833_2071.n291 17.0005
R966 w_833_2071.n299 w_833_2071.n266 17.0005
R967 w_833_2071.n299 w_833_2071.t9 17.0005
R968 w_833_2071.n299 w_833_2071.n265 17.0005
R969 w_833_2071.n299 w_833_2071.n292 17.0005
R970 w_833_2071.n299 w_833_2071.n264 17.0005
R971 w_833_2071.n299 w_833_2071.n293 17.0005
R972 w_833_2071.n299 w_833_2071.n263 17.0005
R973 w_833_2071.n299 w_833_2071.n294 17.0005
R974 w_833_2071.n299 w_833_2071.n262 17.0005
R975 w_833_2071.n299 w_833_2071.n295 17.0005
R976 w_833_2071.n299 w_833_2071.n261 17.0005
R977 w_833_2071.n299 w_833_2071.n296 17.0005
R978 w_833_2071.n299 w_833_2071.n260 17.0005
R979 w_833_2071.n299 w_833_2071.n297 17.0005
R980 w_833_2071.n299 w_833_2071.n259 17.0005
R981 w_833_2071.n299 w_833_2071.n298 17.0005
R982 w_833_2071.n71 w_833_2071.n29 17.0005
R983 w_833_2071.n71 w_833_2071.n30 17.0005
R984 w_833_2071.n71 w_833_2071.n28 17.0005
R985 w_833_2071.n71 w_833_2071.n31 17.0005
R986 w_833_2071.n71 w_833_2071.n27 17.0005
R987 w_833_2071.n71 w_833_2071.n34 17.0005
R988 w_833_2071.n71 w_833_2071.n26 17.0005
R989 w_833_2071.n71 w_833_2071.n35 17.0005
R990 w_833_2071.n71 w_833_2071.n25 17.0005
R991 w_833_2071.n71 w_833_2071.n36 17.0005
R992 w_833_2071.n71 w_833_2071.n23 17.0005
R993 w_833_2071.n71 w_833_2071.n37 17.0005
R994 w_833_2071.n71 w_833_2071.n22 17.0005
R995 w_833_2071.n71 w_833_2071.n38 17.0005
R996 w_833_2071.n71 w_833_2071.n21 17.0005
R997 w_833_2071.n71 w_833_2071.n41 17.0005
R998 w_833_2071.n71 w_833_2071.n20 17.0005
R999 w_833_2071.n71 w_833_2071.n42 17.0005
R1000 w_833_2071.n71 w_833_2071.n19 17.0005
R1001 w_833_2071.n71 w_833_2071.n43 17.0005
R1002 w_833_2071.n71 w_833_2071.n18 17.0005
R1003 w_833_2071.n71 w_833_2071.n44 17.0005
R1004 w_833_2071.n71 w_833_2071.n17 17.0005
R1005 w_833_2071.n71 w_833_2071.n45 17.0005
R1006 w_833_2071.n71 w_833_2071.n16 17.0005
R1007 w_833_2071.n71 w_833_2071.n46 17.0005
R1008 w_833_2071.n71 w_833_2071.n15 17.0005
R1009 w_833_2071.n71 w_833_2071.n47 17.0005
R1010 w_833_2071.n71 w_833_2071.n14 17.0005
R1011 w_833_2071.n71 w_833_2071.n48 17.0005
R1012 w_833_2071.n71 w_833_2071.n10 17.0005
R1013 w_833_2071.n71 w_833_2071.n49 17.0005
R1014 w_833_2071.n71 w_833_2071.n9 17.0005
R1015 w_833_2071.n71 w_833_2071.n50 17.0005
R1016 w_833_2071.n71 w_833_2071.n8 17.0005
R1017 w_833_2071.n71 w_833_2071.n51 17.0005
R1018 w_833_2071.n71 w_833_2071.n6 17.0005
R1019 w_833_2071.n71 w_833_2071.n52 17.0005
R1020 w_833_2071.n71 w_833_2071.n5 17.0005
R1021 w_833_2071.n71 w_833_2071.n53 17.0005
R1022 w_833_2071.n71 w_833_2071.t33 17.0005
R1023 w_833_2071.n322 w_833_2071.n71 17.0005
R1024 w_833_2071.n167 w_833_2071.t124 15.3683
R1025 w_833_2071.n131 w_833_2071.t125 15.3683
R1026 w_833_2071.n295 w_833_2071.t7 15.0475
R1027 w_833_2071.n244 w_833_2071.t83 15.0005
R1028 w_833_2071.n246 w_833_2071.t70 15.0005
R1029 w_833_2071.n247 w_833_2071.t96 15.0005
R1030 w_833_2071.n249 w_833_2071.t92 15.0005
R1031 w_833_2071.n251 w_833_2071.t108 15.0005
R1032 w_833_2071.n253 w_833_2071.t54 15.0005
R1033 w_833_2071.n255 w_833_2071.t72 15.0005
R1034 w_833_2071.n257 w_833_2071.t85 15.0005
R1035 w_833_2071.n315 w_833_2071.t74 15.0005
R1036 w_833_2071.n313 w_833_2071.t100 15.0005
R1037 w_833_2071.n311 w_833_2071.t56 15.0005
R1038 w_833_2071.n309 w_833_2071.t110 15.0005
R1039 w_833_2071.n307 w_833_2071.t58 15.0005
R1040 w_833_2071.n305 w_833_2071.t112 15.0005
R1041 w_833_2071.n303 w_833_2071.t87 15.0005
R1042 w_833_2071.n242 w_833_2071.t68 15.0005
R1043 w_833_2071.n165 w_833_2071.t60 15.0005
R1044 w_833_2071.n163 w_833_2071.t76 15.0005
R1045 w_833_2071.n161 w_833_2071.t64 15.0005
R1046 w_833_2071.n160 w_833_2071.t94 15.0005
R1047 w_833_2071.n158 w_833_2071.t90 15.0005
R1048 w_833_2071.n156 w_833_2071.t102 15.0005
R1049 w_833_2071.n154 w_833_2071.t116 15.0005
R1050 w_833_2071.n152 w_833_2071.t62 15.0005
R1051 w_833_2071.n150 w_833_2071.t78 15.0005
R1052 w_833_2071.n148 w_833_2071.t66 15.0005
R1053 w_833_2071.n146 w_833_2071.t98 15.0005
R1054 w_833_2071.n144 w_833_2071.t114 15.0005
R1055 w_833_2071.n142 w_833_2071.t104 15.0005
R1056 w_833_2071.n140 w_833_2071.t118 15.0005
R1057 w_833_2071.n138 w_833_2071.t106 15.0005
R1058 w_833_2071.n136 w_833_2071.t80 15.0005
R1059 w_833_2071.n167 w_833_2071.t122 14.6976
R1060 w_833_2071.n131 w_833_2071.t123 14.6976
R1061 w_833_2071.n322 w_833_2071.n56 14.1283
R1062 w_833_2071.n258 w_833_2071.n1 13.8647
R1063 w_833_2071.n327 w_833_2071.n326 13.5377
R1064 w_833_2071.n82 w_833_2071.n2 13.5377
R1065 w_833_2071.n190 w_833_2071.n189 13.5377
R1066 w_833_2071.n329 w_833_2071.n328 13.5377
R1067 w_833_2071.n216 w_833_2071.n1 13.5005
R1068 w_833_2071.n188 w_833_2071.n187 13.5005
R1069 w_833_2071.t11 w_833_2071.n51 11.2858
R1070 w_833_2071.n268 w_833_2071.t12 11.2858
R1071 w_833_2071.t18 w_833_2071.n27 11.2858
R1072 w_833_2071.n133 w_833_2071.n132 9.0005
R1073 w_833_2071.n175 w_833_2071.n100 9.0005
R1074 w_833_2071.n169 w_833_2071.n168 9.0005
R1075 w_833_2071.n130 w_833_2071.n89 8.46995
R1076 w_833_2071.n122 w_833_2071.n89 8.46995
R1077 w_833_2071.n172 w_833_2071.n89 8.46995
R1078 w_833_2071.n182 w_833_2071.n89 8.46995
R1079 w_833_2071.n178 w_833_2071.n89 8.46995
R1080 w_833_2071.n116 w_833_2071.n89 8.46995
R1081 w_833_2071.n321 w_833_2071.n207 8.46995
R1082 w_833_2071.n321 w_833_2071.n203 8.46995
R1083 w_833_2071.n321 w_833_2071.n201 8.46995
R1084 w_833_2071.n321 w_833_2071.n210 8.46995
R1085 w_833_2071.n321 w_833_2071.n199 8.46995
R1086 w_833_2071.n321 w_833_2071.n197 8.46995
R1087 w_833_2071.n126 w_833_2071.n89 8.46995
R1088 w_833_2071.t55 w_833_2071.n215 8.46336
R1089 w_833_2071.t61 w_833_2071.n101 8.45649
R1090 w_833_2071.n279 w_833_2071.n53 7.52401
R1091 w_833_2071.n280 w_833_2071.n5 7.52401
R1092 w_833_2071.n278 w_833_2071.n52 7.52401
R1093 w_833_2071.n281 w_833_2071.n6 7.52401
R1094 w_833_2071.n277 w_833_2071.n51 7.52401
R1095 w_833_2071.n282 w_833_2071.n8 7.52401
R1096 w_833_2071.n276 w_833_2071.n50 7.52401
R1097 w_833_2071.n283 w_833_2071.t14 7.52401
R1098 w_833_2071.n283 w_833_2071.n9 7.52401
R1099 w_833_2071.n275 w_833_2071.n49 7.52401
R1100 w_833_2071.n284 w_833_2071.n10 7.52401
R1101 w_833_2071.n274 w_833_2071.n48 7.52401
R1102 w_833_2071.n285 w_833_2071.n14 7.52401
R1103 w_833_2071.n286 w_833_2071.n15 7.52401
R1104 w_833_2071.n272 w_833_2071.n46 7.52401
R1105 w_833_2071.n287 w_833_2071.n16 7.52401
R1106 w_833_2071.n271 w_833_2071.n45 7.52401
R1107 w_833_2071.n288 w_833_2071.n17 7.52401
R1108 w_833_2071.t0 w_833_2071.n17 7.52401
R1109 w_833_2071.n269 w_833_2071.n44 7.52401
R1110 w_833_2071.n289 w_833_2071.n18 7.52401
R1111 w_833_2071.n268 w_833_2071.n43 7.52401
R1112 w_833_2071.n290 w_833_2071.n19 7.52401
R1113 w_833_2071.n267 w_833_2071.n42 7.52401
R1114 w_833_2071.n291 w_833_2071.n20 7.52401
R1115 w_833_2071.n266 w_833_2071.n41 7.52401
R1116 w_833_2071.t9 w_833_2071.n21 7.52401
R1117 w_833_2071.n265 w_833_2071.n38 7.52401
R1118 w_833_2071.n292 w_833_2071.n22 7.52401
R1119 w_833_2071.n264 w_833_2071.n37 7.52401
R1120 w_833_2071.n293 w_833_2071.n23 7.52401
R1121 w_833_2071.n263 w_833_2071.n36 7.52401
R1122 w_833_2071.n294 w_833_2071.n25 7.52401
R1123 w_833_2071.n262 w_833_2071.n35 7.52401
R1124 w_833_2071.n295 w_833_2071.n26 7.52401
R1125 w_833_2071.n261 w_833_2071.n34 7.52401
R1126 w_833_2071.n296 w_833_2071.n27 7.52401
R1127 w_833_2071.n260 w_833_2071.n31 7.52401
R1128 w_833_2071.n297 w_833_2071.n28 7.52401
R1129 w_833_2071.n259 w_833_2071.t81 7.52401
R1130 w_833_2071.n259 w_833_2071.n30 7.52401
R1131 w_833_2071.n298 w_833_2071.n29 7.52401
R1132 w_833_2071.n33 w_833_2071.t127 6.43891
R1133 w_833_2071.n78 w_833_2071.t129 6.43891
R1134 w_833_2071.n96 w_833_2071.t140 6.43891
R1135 w_833_2071.n63 w_833_2071.t136 6.43891
R1136 w_833_2071.n55 w_833_2071.t146 6.4061
R1137 w_833_2071.n87 w_833_2071.t139 6.4061
R1138 w_833_2071.n195 w_833_2071.t34 6.4061
R1139 w_833_2071.n70 w_833_2071.t42 6.4061
R1140 w_833_2071.n168 w_833_2071.n167 6.15663
R1141 w_833_2071.n132 w_833_2071.n131 6.15663
R1142 w_833_2071.n54 w_833_2071.t6 6.12323
R1143 w_833_2071.n12 w_833_2071.t47 6.12323
R1144 w_833_2071.n11 w_833_2071.t4 6.12323
R1145 w_833_2071.n4 w_833_2071.t35 6.12323
R1146 w_833_2071.n39 w_833_2071.t36 6.12323
R1147 w_833_2071.n32 w_833_2071.t19 6.12323
R1148 w_833_2071.n86 w_833_2071.t48 6.12323
R1149 w_833_2071.n73 w_833_2071.t21 6.12323
R1150 w_833_2071.n84 w_833_2071.t3 6.12323
R1151 w_833_2071.n80 w_833_2071.t31 6.12323
R1152 w_833_2071.n79 w_833_2071.t126 6.12323
R1153 w_833_2071.n77 w_833_2071.t25 6.12323
R1154 w_833_2071.n194 w_833_2071.t30 6.12323
R1155 w_833_2071.n91 w_833_2071.t15 6.12323
R1156 w_833_2071.n192 w_833_2071.t40 6.12323
R1157 w_833_2071.n98 w_833_2071.t24 6.12323
R1158 w_833_2071.n97 w_833_2071.t17 6.12323
R1159 w_833_2071.n95 w_833_2071.t22 6.12323
R1160 w_833_2071.t55 w_833_2071.n227 6.12323
R1161 w_833_2071.n69 w_833_2071.t45 6.12323
R1162 w_833_2071.n58 w_833_2071.t53 6.12323
R1163 w_833_2071.n67 w_833_2071.t44 6.12323
R1164 w_833_2071.n65 w_833_2071.t10 6.12323
R1165 w_833_2071.n64 w_833_2071.t28 6.12323
R1166 w_833_2071.n62 w_833_2071.t8 6.12323
R1167 w_833_2071.t61 w_833_2071.n185 6.12223
R1168 w_833_2071.n326 w_833_2071.t13 5.67005
R1169 w_833_2071.n82 w_833_2071.t26 5.67005
R1170 w_833_2071.n190 w_833_2071.t49 5.67005
R1171 w_833_2071.t1 w_833_2071.n329 5.67005
R1172 w_833_2071.n170 w_833_2071.n89 5.61281
R1173 w_833_2071.n174 w_833_2071.n89 5.61281
R1174 w_833_2071.n184 w_833_2071.n89 5.61281
R1175 w_833_2071.n180 w_833_2071.n89 5.61281
R1176 w_833_2071.n176 w_833_2071.n89 5.61281
R1177 w_833_2071.n321 w_833_2071.n205 5.61281
R1178 w_833_2071.n321 w_833_2071.n204 5.61281
R1179 w_833_2071.n321 w_833_2071.n208 5.61281
R1180 w_833_2071.n321 w_833_2071.n202 5.61281
R1181 w_833_2071.n321 w_833_2071.n209 5.61281
R1182 w_833_2071.n321 w_833_2071.n200 5.61281
R1183 w_833_2071.n321 w_833_2071.n211 5.61281
R1184 w_833_2071.n321 w_833_2071.n198 5.61281
R1185 w_833_2071.n321 w_833_2071.n320 5.61281
R1186 w_833_2071.n124 w_833_2071.n89 5.61281
R1187 w_833_2071.n120 w_833_2071.n89 5.61281
R1188 w_833_2071.n118 w_833_2071.n89 5.61281
R1189 w_833_2071.n128 w_833_2071.n89 5.61121
R1190 w_833_2071.n321 w_833_2071.n206 5.61121
R1191 w_833_2071.t61 w_833_2071.n113 5.56245
R1192 w_833_2071.t61 w_833_2071.n112 5.56245
R1193 w_833_2071.t61 w_833_2071.n111 5.56245
R1194 w_833_2071.t61 w_833_2071.n110 5.56245
R1195 w_833_2071.t61 w_833_2071.n109 5.56245
R1196 w_833_2071.t61 w_833_2071.n108 5.56245
R1197 w_833_2071.t61 w_833_2071.n107 5.56245
R1198 w_833_2071.t55 w_833_2071.n318 5.56245
R1199 w_833_2071.n319 w_833_2071.t55 5.56245
R1200 w_833_2071.t55 w_833_2071.n229 5.56245
R1201 w_833_2071.t55 w_833_2071.n226 5.56245
R1202 w_833_2071.t55 w_833_2071.n224 5.56245
R1203 w_833_2071.t55 w_833_2071.n222 5.56245
R1204 w_833_2071.t55 w_833_2071.n220 5.56245
R1205 w_833_2071.t55 w_833_2071.n231 5.56245
R1206 w_833_2071.t55 w_833_2071.n233 5.56245
R1207 w_833_2071.t55 w_833_2071.n235 5.56245
R1208 w_833_2071.t55 w_833_2071.n237 5.56245
R1209 w_833_2071.t55 w_833_2071.n239 5.56245
R1210 w_833_2071.t55 w_833_2071.n241 5.56245
R1211 w_833_2071.n301 w_833_2071.t89 5.56245
R1212 w_833_2071.t55 w_833_2071.n214 5.56245
R1213 w_833_2071.t61 w_833_2071.n106 5.56245
R1214 w_833_2071.t61 w_833_2071.n105 5.56245
R1215 w_833_2071.t61 w_833_2071.n104 5.56245
R1216 w_833_2071.t61 w_833_2071.n103 5.56245
R1217 w_833_2071.t61 w_833_2071.n114 5.56245
R1218 w_833_2071.t61 w_833_2071.n115 5.56245
R1219 w_833_2071.t61 w_833_2071.n166 5.56245
R1220 w_833_2071.n135 w_833_2071.t82 5.56245
R1221 w_833_2071.n188 w_833_2071.n100 4.72356
R1222 w_833_2071.n299 w_833_2071.n56 4.25726
R1223 w_833_2071.n273 w_833_2071.t43 3.76226
R1224 w_833_2071.t43 w_833_2071.n47 3.76226
R1225 w_833_2071.t16 w_833_2071.n36 3.76226
R1226 w_833_2071.n196 w_833_2071.n94 3.30365
R1227 w_833_2071.n196 w_833_2071.n99 3.30365
R1228 w_833_2071.n196 w_833_2071.n93 3.30365
R1229 w_833_2071.n196 w_833_2071.n193 3.30365
R1230 w_833_2071.n196 w_833_2071.n92 3.30365
R1231 w_833_2071.n196 w_833_2071.n195 3.30365
R1232 w_833_2071.n88 w_833_2071.n76 3.30365
R1233 w_833_2071.n88 w_833_2071.n81 3.30365
R1234 w_833_2071.n88 w_833_2071.n75 3.30365
R1235 w_833_2071.n88 w_833_2071.n85 3.30365
R1236 w_833_2071.n88 w_833_2071.n74 3.30365
R1237 w_833_2071.n88 w_833_2071.n87 3.30365
R1238 w_833_2071.n323 w_833_2071.n24 3.30365
R1239 w_833_2071.n323 w_833_2071.n40 3.30365
R1240 w_833_2071.n324 w_833_2071.n323 3.30365
R1241 w_833_2071.n323 w_833_2071.n3 3.30365
R1242 w_833_2071.n323 w_833_2071.n13 3.30365
R1243 w_833_2071.n323 w_833_2071.n55 3.30365
R1244 w_833_2071.n71 w_833_2071.n61 3.30365
R1245 w_833_2071.n71 w_833_2071.n66 3.30365
R1246 w_833_2071.n71 w_833_2071.n60 3.30365
R1247 w_833_2071.n71 w_833_2071.n68 3.30365
R1248 w_833_2071.n71 w_833_2071.n59 3.30365
R1249 w_833_2071.n71 w_833_2071.n70 3.30365
R1250 w_833_2071.n196 w_833_2071.n90 2.71714
R1251 w_833_2071.n88 w_833_2071.n72 2.71714
R1252 w_833_2071.n323 w_833_2071.n7 2.71714
R1253 w_833_2071.n71 w_833_2071.n57 2.71714
R1254 w_833_2071.n196 w_833_2071.n96 2.71618
R1255 w_833_2071.n88 w_833_2071.n78 2.71618
R1256 w_833_2071.n323 w_833_2071.n33 2.71618
R1257 w_833_2071.n71 w_833_2071.n63 2.71618
R1258 w_833_2071.n168 w_833_2071.n100 2.10491
R1259 w_833_2071.n132 w_833_2071.n100 2.10491
R1260 w_833_2071.n270 w_833_2071.n213 1.14089
R1261 w_833_2071.n302 w_833_2071.n300 1.13323
R1262 w_833_2071.n300 w_833_2071.n258 1.05833
R1263 w_833_2071.n270 w_833_2071.n258 1.04625
R1264 w_833_2071.n328 w_833_2071.n1 0.80919
R1265 w_833_2071.n166 w_833_2071.n165 0.80612
R1266 w_833_2071.n136 w_833_2071.n135 0.805774
R1267 w_833_2071.n189 w_833_2071.n2 0.794017
R1268 w_833_2071.n328 w_833_2071.n327 0.789466
R1269 w_833_2071.n327 w_833_2071.n2 0.789466
R1270 w_833_2071.n320 w_833_2071.n319 0.722964
R1271 w_833_2071.n301 w_833_2071.n205 0.693971
R1272 w_833_2071.n189 w_833_2071.n188 0.693879
R1273 w_833_2071.n247 w_833_2071.n246 0.6055
R1274 w_833_2071.n161 w_833_2071.n160 0.6055
R1275 w_833_2071.n169 w_833_2071.n166 0.596545
R1276 w_833_2071.n135 w_833_2071.n134 0.569391
R1277 w_833_2071.n241 w_833_2071.n240 0.562058
R1278 w_833_2071.n177 w_833_2071.n106 0.562058
R1279 w_833_2071.n179 w_833_2071.n105 0.562058
R1280 w_833_2071.n181 w_833_2071.n104 0.562058
R1281 w_833_2071.n183 w_833_2071.n103 0.562058
R1282 w_833_2071.n173 w_833_2071.n114 0.562058
R1283 w_833_2071.n171 w_833_2071.n115 0.562058
R1284 w_833_2071.n129 w_833_2071.n113 0.561712
R1285 w_833_2071.n127 w_833_2071.n112 0.561712
R1286 w_833_2071.n125 w_833_2071.n111 0.561712
R1287 w_833_2071.n123 w_833_2071.n110 0.561712
R1288 w_833_2071.n121 w_833_2071.n109 0.561712
R1289 w_833_2071.n119 w_833_2071.n108 0.561712
R1290 w_833_2071.n117 w_833_2071.n107 0.561712
R1291 w_833_2071.n318 w_833_2071.n317 0.561712
R1292 w_833_2071.n229 w_833_2071.n228 0.561712
R1293 w_833_2071.n226 w_833_2071.n225 0.561712
R1294 w_833_2071.n224 w_833_2071.n223 0.561712
R1295 w_833_2071.n222 w_833_2071.n221 0.561712
R1296 w_833_2071.n220 w_833_2071.n219 0.561712
R1297 w_833_2071.n231 w_833_2071.n230 0.561712
R1298 w_833_2071.n233 w_833_2071.n232 0.561712
R1299 w_833_2071.n235 w_833_2071.n234 0.561712
R1300 w_833_2071.n237 w_833_2071.n236 0.561712
R1301 w_833_2071.n239 w_833_2071.n238 0.561712
R1302 w_833_2071.n214 w_833_2071.n212 0.561712
R1303 w_833_2071.n137 w_833_2071.n113 0.50362
R1304 w_833_2071.n139 w_833_2071.n112 0.50362
R1305 w_833_2071.n141 w_833_2071.n111 0.50362
R1306 w_833_2071.n143 w_833_2071.n110 0.50362
R1307 w_833_2071.n145 w_833_2071.n109 0.50362
R1308 w_833_2071.n147 w_833_2071.n108 0.50362
R1309 w_833_2071.n149 w_833_2071.n107 0.50362
R1310 w_833_2071.n318 w_833_2071.n316 0.50362
R1311 w_833_2071.n319 w_833_2071.n213 0.50362
R1312 w_833_2071.n245 w_833_2071.n229 0.50362
R1313 w_833_2071.n248 w_833_2071.n226 0.50362
R1314 w_833_2071.n250 w_833_2071.n224 0.50362
R1315 w_833_2071.n252 w_833_2071.n222 0.50362
R1316 w_833_2071.n254 w_833_2071.n220 0.50362
R1317 w_833_2071.n314 w_833_2071.n231 0.50362
R1318 w_833_2071.n312 w_833_2071.n233 0.50362
R1319 w_833_2071.n310 w_833_2071.n235 0.50362
R1320 w_833_2071.n308 w_833_2071.n237 0.50362
R1321 w_833_2071.n306 w_833_2071.n239 0.50362
R1322 w_833_2071.n302 w_833_2071.n301 0.50362
R1323 w_833_2071.n243 w_833_2071.n214 0.50362
R1324 w_833_2071.n304 w_833_2071.n241 0.503274
R1325 w_833_2071.n153 w_833_2071.n106 0.503274
R1326 w_833_2071.n155 w_833_2071.n105 0.503274
R1327 w_833_2071.n157 w_833_2071.n104 0.503274
R1328 w_833_2071.n159 w_833_2071.n103 0.503274
R1329 w_833_2071.n162 w_833_2071.n114 0.503274
R1330 w_833_2071.n164 w_833_2071.n115 0.503274
R1331 w_833_2071.n299 w_833_2071.n270 0.499574
R1332 w_833_2071.n300 w_833_2071.n299 0.498883
R1333 w_833_2071.n326 w_833_2071.n325 0.37848
R1334 w_833_2071.n83 w_833_2071.n82 0.37848
R1335 w_833_2071.n191 w_833_2071.n190 0.37848
R1336 w_833_2071.n329 w_833_2071.n0 0.37848
R1337 w_833_2071.n32 w_833_2071.n24 0.365272
R1338 w_833_2071.n77 w_833_2071.n76 0.365272
R1339 w_833_2071.n95 w_833_2071.n94 0.365272
R1340 w_833_2071.n62 w_833_2071.n61 0.365272
R1341 w_833_2071.n13 w_833_2071.n12 0.364033
R1342 w_833_2071.n74 w_833_2071.n73 0.364033
R1343 w_833_2071.n92 w_833_2071.n91 0.364033
R1344 w_833_2071.n59 w_833_2071.n58 0.364033
R1345 w_833_2071.n55 w_833_2071.n54 0.357939
R1346 w_833_2071.n87 w_833_2071.n86 0.357939
R1347 w_833_2071.n195 w_833_2071.n194 0.357939
R1348 w_833_2071.n70 w_833_2071.n69 0.357939
R1349 w_833_2071.n151 w_833_2071.n101 0.354712
R1350 w_833_2071.n40 w_833_2071.n39 0.343272
R1351 w_833_2071.n81 w_833_2071.n79 0.343272
R1352 w_833_2071.n99 w_833_2071.n97 0.343272
R1353 w_833_2071.n66 w_833_2071.n64 0.343272
R1354 w_833_2071.n11 w_833_2071.n3 0.342033
R1355 w_833_2071.n85 w_833_2071.n84 0.342033
R1356 w_833_2071.n193 w_833_2071.n192 0.342033
R1357 w_833_2071.n68 w_833_2071.n67 0.342033
R1358 w_833_2071.n256 w_833_2071.n215 0.340978
R1359 w_833_2071.n324 w_833_2071.n4 0.321272
R1360 w_833_2071.n80 w_833_2071.n75 0.321272
R1361 w_833_2071.n98 w_833_2071.n93 0.321272
R1362 w_833_2071.n65 w_833_2071.n60 0.321272
R1363 w_833_2071.n54 w_833_2071.n7 0.320626
R1364 w_833_2071.n86 w_833_2071.n72 0.320626
R1365 w_833_2071.n194 w_833_2071.n90 0.320626
R1366 w_833_2071.n69 w_833_2071.n57 0.320626
R1367 w_833_2071.n325 w_833_2071.n324 0.320033
R1368 w_833_2071.n83 w_833_2071.n75 0.320033
R1369 w_833_2071.n191 w_833_2071.n93 0.320033
R1370 w_833_2071.n60 w_833_2071.n0 0.320033
R1371 w_833_2071.n33 w_833_2071.n32 0.319212
R1372 w_833_2071.n78 w_833_2071.n77 0.319212
R1373 w_833_2071.n96 w_833_2071.n95 0.319212
R1374 w_833_2071.n63 w_833_2071.n62 0.319212
R1375 w_833_2071.n12 w_833_2071.n7 0.315027
R1376 w_833_2071.n73 w_833_2071.n72 0.315027
R1377 w_833_2071.n91 w_833_2071.n90 0.315027
R1378 w_833_2071.n58 w_833_2071.n57 0.315027
R1379 w_833_2071.n218 w_833_2071.n217 0.305134
R1380 w_833_2071.n242 w_833_2071.n213 0.303
R1381 w_833_2071.n243 w_833_2071.n242 0.303
R1382 w_833_2071.n244 w_833_2071.n243 0.303
R1383 w_833_2071.n245 w_833_2071.n244 0.303
R1384 w_833_2071.n246 w_833_2071.n245 0.303
R1385 w_833_2071.n248 w_833_2071.n247 0.303
R1386 w_833_2071.n249 w_833_2071.n248 0.303
R1387 w_833_2071.n250 w_833_2071.n249 0.303
R1388 w_833_2071.n251 w_833_2071.n250 0.303
R1389 w_833_2071.n252 w_833_2071.n251 0.303
R1390 w_833_2071.n253 w_833_2071.n252 0.303
R1391 w_833_2071.n254 w_833_2071.n253 0.303
R1392 w_833_2071.n255 w_833_2071.n254 0.303
R1393 w_833_2071.n256 w_833_2071.n255 0.303
R1394 w_833_2071.n257 w_833_2071.n256 0.303
R1395 w_833_2071.n316 w_833_2071.n257 0.303
R1396 w_833_2071.n316 w_833_2071.n315 0.303
R1397 w_833_2071.n315 w_833_2071.n314 0.303
R1398 w_833_2071.n314 w_833_2071.n313 0.303
R1399 w_833_2071.n313 w_833_2071.n312 0.303
R1400 w_833_2071.n312 w_833_2071.n311 0.303
R1401 w_833_2071.n311 w_833_2071.n310 0.303
R1402 w_833_2071.n310 w_833_2071.n309 0.303
R1403 w_833_2071.n309 w_833_2071.n308 0.303
R1404 w_833_2071.n308 w_833_2071.n307 0.303
R1405 w_833_2071.n307 w_833_2071.n306 0.303
R1406 w_833_2071.n306 w_833_2071.n305 0.303
R1407 w_833_2071.n305 w_833_2071.n304 0.303
R1408 w_833_2071.n304 w_833_2071.n303 0.303
R1409 w_833_2071.n303 w_833_2071.n302 0.303
R1410 w_833_2071.n165 w_833_2071.n164 0.303
R1411 w_833_2071.n164 w_833_2071.n163 0.303
R1412 w_833_2071.n163 w_833_2071.n162 0.303
R1413 w_833_2071.n162 w_833_2071.n161 0.303
R1414 w_833_2071.n160 w_833_2071.n159 0.303
R1415 w_833_2071.n159 w_833_2071.n158 0.303
R1416 w_833_2071.n158 w_833_2071.n157 0.303
R1417 w_833_2071.n157 w_833_2071.n156 0.303
R1418 w_833_2071.n156 w_833_2071.n155 0.303
R1419 w_833_2071.n155 w_833_2071.n154 0.303
R1420 w_833_2071.n154 w_833_2071.n153 0.303
R1421 w_833_2071.n153 w_833_2071.n152 0.303
R1422 w_833_2071.n152 w_833_2071.n151 0.303
R1423 w_833_2071.n151 w_833_2071.n150 0.303
R1424 w_833_2071.n150 w_833_2071.n149 0.303
R1425 w_833_2071.n149 w_833_2071.n148 0.303
R1426 w_833_2071.n148 w_833_2071.n147 0.303
R1427 w_833_2071.n147 w_833_2071.n146 0.303
R1428 w_833_2071.n146 w_833_2071.n145 0.303
R1429 w_833_2071.n145 w_833_2071.n144 0.303
R1430 w_833_2071.n144 w_833_2071.n143 0.303
R1431 w_833_2071.n143 w_833_2071.n142 0.303
R1432 w_833_2071.n142 w_833_2071.n141 0.303
R1433 w_833_2071.n141 w_833_2071.n140 0.303
R1434 w_833_2071.n140 w_833_2071.n139 0.303
R1435 w_833_2071.n139 w_833_2071.n138 0.303
R1436 w_833_2071.n138 w_833_2071.n137 0.303
R1437 w_833_2071.n137 w_833_2071.n136 0.303
R1438 w_833_2071.n325 w_833_2071.n3 0.299272
R1439 w_833_2071.n85 w_833_2071.n83 0.299272
R1440 w_833_2071.n193 w_833_2071.n191 0.299272
R1441 w_833_2071.n68 w_833_2071.n0 0.299272
R1442 w_833_2071.n40 w_833_2071.n4 0.298033
R1443 w_833_2071.n81 w_833_2071.n80 0.298033
R1444 w_833_2071.n99 w_833_2071.n98 0.298033
R1445 w_833_2071.n66 w_833_2071.n65 0.298033
R1446 w_833_2071.n186 w_833_2071.n102 0.277397
R1447 w_833_2071.n13 w_833_2071.n11 0.277272
R1448 w_833_2071.n84 w_833_2071.n74 0.277272
R1449 w_833_2071.n192 w_833_2071.n92 0.277272
R1450 w_833_2071.n67 w_833_2071.n59 0.277272
R1451 w_833_2071.n39 w_833_2071.n24 0.276033
R1452 w_833_2071.n79 w_833_2071.n76 0.276033
R1453 w_833_2071.n97 w_833_2071.n94 0.276033
R1454 w_833_2071.n64 w_833_2071.n61 0.276033
R1455 w_833_2071.n230 w_833_2071.n202 0.198759
R1456 w_833_2071.n119 w_833_2071.n118 0.198419
R1457 w_833_2071.n185 w_833_2071.n184 0.191425
R1458 w_833_2071.n227 w_833_2071.n211 0.191086
R1459 w_833_2071.n240 w_833_2071.n205 0.191086
R1460 w_833_2071.n317 w_833_2071.n201 0.187772
R1461 w_833_2071.n117 w_833_2071.n116 0.187772
R1462 w_833_2071.n240 w_833_2071.n206 0.186494
R1463 w_833_2071.n129 w_833_2071.n128 0.186494
R1464 w_833_2071.n227 w_833_2071.n198 0.184092
R1465 w_833_2071.n185 w_833_2071.n174 0.183752
R1466 w_833_2071.n225 w_833_2071.n199 0.180439
R1467 w_833_2071.n238 w_833_2071.n207 0.180439
R1468 w_833_2071.n183 w_833_2071.n182 0.180439
R1469 w_833_2071.n127 w_833_2071.n126 0.180439
R1470 w_833_2071.n217 w_833_2071.n209 0.176759
R1471 w_833_2071.n230 w_833_2071.n208 0.176419
R1472 w_833_2071.n120 w_833_2071.n119 0.176419
R1473 w_833_2071.n228 w_833_2071.n197 0.173106
R1474 w_833_2071.n173 w_833_2071.n172 0.173106
R1475 w_833_2071.n176 w_833_2071.n175 0.172752
R1476 w_833_2071.n236 w_833_2071.n204 0.169425
R1477 w_833_2071.n181 w_833_2071.n180 0.169425
R1478 w_833_2071.n223 w_833_2071.n200 0.169086
R1479 w_833_2071.n125 w_833_2071.n124 0.169086
R1480 w_833_2071.n219 w_833_2071.n210 0.165772
R1481 w_833_2071.n232 w_833_2071.n203 0.165772
R1482 w_833_2071.n178 w_833_2071.n177 0.165772
R1483 w_833_2071.n122 w_833_2071.n121 0.165772
R1484 w_833_2071.n320 w_833_2071.n212 0.162092
R1485 w_833_2071.n171 w_833_2071.n170 0.161752
R1486 w_833_2071.n221 w_833_2071.n210 0.158439
R1487 w_833_2071.n234 w_833_2071.n203 0.158439
R1488 w_833_2071.n179 w_833_2071.n178 0.158439
R1489 w_833_2071.n123 w_833_2071.n122 0.158439
R1490 w_833_2071.n221 w_833_2071.n200 0.154759
R1491 w_833_2071.n124 w_833_2071.n123 0.154759
R1492 w_833_2071.n234 w_833_2071.n204 0.154419
R1493 w_833_2071.n180 w_833_2071.n179 0.154419
R1494 w_833_2071.n133 w_833_2071.n130 0.152939
R1495 w_833_2071.n212 w_833_2071.n197 0.151106
R1496 w_833_2071.n172 w_833_2071.n171 0.151106
R1497 w_833_2071.n232 w_833_2071.n208 0.147425
R1498 w_833_2071.n177 w_833_2071.n176 0.147425
R1499 w_833_2071.n121 w_833_2071.n120 0.147425
R1500 w_833_2071.n219 w_833_2071.n209 0.147086
R1501 w_833_2071.n187 w_833_2071.n101 0.146921
R1502 w_833_2071.n223 w_833_2071.n199 0.143772
R1503 w_833_2071.n236 w_833_2071.n207 0.143772
R1504 w_833_2071.n182 w_833_2071.n181 0.143772
R1505 w_833_2071.n126 w_833_2071.n125 0.143772
R1506 w_833_2071.n174 w_833_2071.n173 0.140092
R1507 w_833_2071.n228 w_833_2071.n198 0.139752
R1508 w_833_2071.n238 w_833_2071.n206 0.137241
R1509 w_833_2071.n128 w_833_2071.n127 0.137241
R1510 w_833_2071.n217 w_833_2071.n201 0.136439
R1511 w_833_2071.n116 w_833_2071.n102 0.136439
R1512 w_833_2071.n225 w_833_2071.n211 0.132759
R1513 w_833_2071.n184 w_833_2071.n183 0.132419
R1514 w_833_2071.n130 w_833_2071.n129 0.129106
R1515 w_833_2071.n170 w_833_2071.n169 0.127259
R1516 w_833_2071.n118 w_833_2071.n117 0.125425
R1517 w_833_2071.n317 w_833_2071.n202 0.125086
R1518 w_833_2071.n218 w_833_2071.n216 0.1105
R1519 w_833_2071.n216 w_833_2071.n215 0.0990487
R1520 w_833_2071.n187 w_833_2071.n186 0.0763621
R1521 w_833_2071.n134 w_833_2071.n133 0.0353333
R1522 w_833_2071.n175 w_833_2071.n102 0.00416667
R1523 vinp.n0 vinp.t16 15.8289
R1524 vinp.n22 vinp.t27 15.8289
R1525 vinp.n15 vinp.t21 15.6055
R1526 vinp.n7 vinp.t12 15.6055
R1527 vinp.n6 vinp.t13 15.2239
R1528 vinp.n5 vinp.t18 15.2239
R1529 vinp.n4 vinp.t24 15.2239
R1530 vinp.n3 vinp.t7 15.2239
R1531 vinp.n2 vinp.t5 15.2239
R1532 vinp.n1 vinp.t14 15.2239
R1533 vinp.n0 vinp.t9 15.2239
R1534 vinp.n28 vinp.t26 15.2239
R1535 vinp.n27 vinp.t31 15.2239
R1536 vinp.n26 vinp.t2 15.2239
R1537 vinp.n25 vinp.t15 15.2239
R1538 vinp.n24 vinp.t10 15.2239
R1539 vinp.n23 vinp.t25 15.2239
R1540 vinp.n22 vinp.t19 15.2239
R1541 vinp.n15 vinp.t28 15.0005
R1542 vinp.n16 vinp.t8 15.0005
R1543 vinp.n17 vinp.t1 15.0005
R1544 vinp.n18 vinp.t4 15.0005
R1545 vinp.n19 vinp.t0 15.0005
R1546 vinp.n20 vinp.t3 15.0005
R1547 vinp.n21 vinp.t20 15.0005
R1548 vinp.n7 vinp.t17 15.0005
R1549 vinp.n8 vinp.t6 15.0005
R1550 vinp.n9 vinp.t23 15.0005
R1551 vinp.n10 vinp.t30 15.0005
R1552 vinp.n11 vinp.t22 15.0005
R1553 vinp.n12 vinp.t29 15.0005
R1554 vinp.n13 vinp.t11 15.0005
R1555 vinp vinp.n30 12.0616
R1556 vinp.n14 vinp 10.4452
R1557 vinp.n29 vinp 10.1782
R1558 vinp.n29 vinp 9.53331
R1559 vinp.n14 vinp 9.26175
R1560 vinp vinp.n6 4.90238
R1561 vinp vinp.n28 4.90238
R1562 vinp.n1 vinp.n0 0.6055
R1563 vinp.n2 vinp.n1 0.6055
R1564 vinp.n3 vinp.n2 0.6055
R1565 vinp.n4 vinp.n3 0.6055
R1566 vinp.n5 vinp.n4 0.6055
R1567 vinp.n6 vinp.n5 0.6055
R1568 vinp.n23 vinp.n22 0.6055
R1569 vinp.n24 vinp.n23 0.6055
R1570 vinp.n25 vinp.n24 0.6055
R1571 vinp.n26 vinp.n25 0.6055
R1572 vinp.n27 vinp.n26 0.6055
R1573 vinp.n28 vinp.n27 0.6055
R1574 vinp.n16 vinp.n15 0.6055
R1575 vinp.n17 vinp.n16 0.6055
R1576 vinp.n18 vinp.n17 0.6055
R1577 vinp.n19 vinp.n18 0.6055
R1578 vinp.n20 vinp.n19 0.6055
R1579 vinp.n21 vinp.n20 0.6055
R1580 vinp.n8 vinp.n7 0.6055
R1581 vinp.n9 vinp.n8 0.6055
R1582 vinp.n10 vinp.n9 0.6055
R1583 vinp.n11 vinp.n10 0.6055
R1584 vinp.n12 vinp.n11 0.6055
R1585 vinp.n13 vinp.n12 0.6055
R1586 vinp.n30 vinp.n29 0.425328
R1587 vinp vinp.n21 0.333938
R1588 vinp vinp.n13 0.333938
R1589 vinp.n30 vinp.n14 0.241741
R1590 a_610_6649.n10 a_610_6649.t22 18.8663
R1591 a_610_6649.n3 a_610_6649.t15 18.8633
R1592 a_610_6649.n14 a_610_6649.t23 18.619
R1593 a_610_6649.n6 a_610_6649.t16 18.619
R1594 a_610_6649.n12 a_610_6649.t14 18.1315
R1595 a_610_6649.n11 a_610_6649.t13 18.1315
R1596 a_610_6649.n10 a_610_6649.t19 18.1315
R1597 a_610_6649.n5 a_610_6649.t20 18.1285
R1598 a_610_6649.n4 a_610_6649.t27 18.1285
R1599 a_610_6649.n3 a_610_6649.t26 18.1285
R1600 a_610_6649.n16 a_610_6649.t21 17.8842
R1601 a_610_6649.n15 a_610_6649.t18 17.8842
R1602 a_610_6649.n14 a_610_6649.t25 17.8842
R1603 a_610_6649.n8 a_610_6649.t12 17.8842
R1604 a_610_6649.n7 a_610_6649.t24 17.8842
R1605 a_610_6649.n6 a_610_6649.t17 17.8842
R1606 a_610_6649.n18 a_610_6649.n17 15.7467
R1607 a_610_6649.n17 a_610_6649.n16 13.4687
R1608 a_610_6649.n9 a_610_6649.n8 13.4687
R1609 a_610_6649.n9 a_610_6649.n5 11.1279
R1610 a_610_6649.n36 a_610_6649.n18 10.8121
R1611 a_610_6649.n13 a_610_6649.n12 10.3711
R1612 a_610_6649.n27 a_610_6649.n18 9.36767
R1613 a_610_6649.n28 a_610_6649.t7 5.63764
R1614 a_610_6649.n35 a_610_6649.t5 5.63764
R1615 a_610_6649.n26 a_610_6649.t3 5.63764
R1616 a_610_6649.t1 a_610_6649.n37 5.63764
R1617 a_610_6649.n37 a_610_6649.n36 5.47532
R1618 a_610_6649.n27 a_610_6649.n26 5.47498
R1619 a_610_6649.n28 a_610_6649.n27 4.57374
R1620 a_610_6649.n36 a_610_6649.n35 4.57374
R1621 a_610_6649.n23 a_610_6649.t34 4.42794
R1622 a_610_6649.n19 a_610_6649.t29 4.42666
R1623 a_610_6649.n0 a_610_6649.t28 4.42666
R1624 a_610_6649.n29 a_610_6649.t35 4.42557
R1625 a_610_6649.n19 a_610_6649.t33 2.82253
R1626 a_610_6649.n20 a_610_6649.t4 2.82253
R1627 a_610_6649.n33 a_610_6649.t10 2.82253
R1628 a_610_6649.n32 a_610_6649.t11 2.82253
R1629 a_610_6649.n30 a_610_6649.t6 2.82253
R1630 a_610_6649.n29 a_610_6649.t31 2.82253
R1631 a_610_6649.n0 a_610_6649.t32 2.82253
R1632 a_610_6649.n1 a_610_6649.t0 2.82253
R1633 a_610_6649.n21 a_610_6649.t8 2.82253
R1634 a_610_6649.n22 a_610_6649.t9 2.82253
R1635 a_610_6649.n24 a_610_6649.t2 2.82253
R1636 a_610_6649.n23 a_610_6649.t30 2.82253
R1637 a_610_6649.n20 a_610_6649.n19 1.60563
R1638 a_610_6649.n33 a_610_6649.n32 1.60563
R1639 a_610_6649.n30 a_610_6649.n29 1.60563
R1640 a_610_6649.n1 a_610_6649.n0 1.60563
R1641 a_610_6649.n22 a_610_6649.n21 1.60563
R1642 a_610_6649.n24 a_610_6649.n23 1.60563
R1643 a_610_6649.n13 a_610_6649.n9 1.4635
R1644 a_610_6649.n34 a_610_6649.n20 0.803704
R1645 a_610_6649.n32 a_610_6649.n31 0.803704
R1646 a_610_6649.n2 a_610_6649.n1 0.803704
R1647 a_610_6649.n25 a_610_6649.n22 0.803704
R1648 a_610_6649.n34 a_610_6649.n33 0.802423
R1649 a_610_6649.n31 a_610_6649.n30 0.802423
R1650 a_610_6649.n21 a_610_6649.n2 0.802423
R1651 a_610_6649.n25 a_610_6649.n24 0.802423
R1652 a_610_6649.n17 a_610_6649.n13 0.7463
R1653 a_610_6649.n15 a_610_6649.n14 0.7353
R1654 a_610_6649.n16 a_610_6649.n15 0.7353
R1655 a_610_6649.n11 a_610_6649.n10 0.7353
R1656 a_610_6649.n12 a_610_6649.n11 0.7353
R1657 a_610_6649.n7 a_610_6649.n6 0.7353
R1658 a_610_6649.n8 a_610_6649.n7 0.7353
R1659 a_610_6649.n4 a_610_6649.n3 0.7353
R1660 a_610_6649.n5 a_610_6649.n4 0.7353
R1661 a_610_6649.n31 a_610_6649.n28 0.390831
R1662 a_610_6649.n35 a_610_6649.n34 0.390831
R1663 a_610_6649.n26 a_610_6649.n25 0.390831
R1664 a_610_6649.n37 a_610_6649.n2 0.390492
R1665 vinn.n15 vinn.t28 15.8289
R1666 vinn.n7 vinn.t18 15.8289
R1667 vinn.n0 vinn.t9 15.6055
R1668 vinn.n22 vinn.t20 15.6055
R1669 vinn.n21 vinn.t26 15.2239
R1670 vinn.n20 vinn.t0 15.2239
R1671 vinn.n19 vinn.t4 15.2239
R1672 vinn.n18 vinn.t13 15.2239
R1673 vinn.n17 vinn.t10 15.2239
R1674 vinn.n16 vinn.t27 15.2239
R1675 vinn.n15 vinn.t21 15.2239
R1676 vinn.n13 vinn.t15 15.2239
R1677 vinn.n12 vinn.t22 15.2239
R1678 vinn.n11 vinn.t29 15.2239
R1679 vinn.n10 vinn.t8 15.2239
R1680 vinn.n9 vinn.t5 15.2239
R1681 vinn.n8 vinn.t14 15.2239
R1682 vinn.n7 vinn.t12 15.2239
R1683 vinn.n0 vinn.t11 15.0005
R1684 vinn.n1 vinn.t2 15.0005
R1685 vinn.n2 vinn.t19 15.0005
R1686 vinn.n3 vinn.t24 15.0005
R1687 vinn.n4 vinn.t16 15.0005
R1688 vinn.n5 vinn.t23 15.0005
R1689 vinn.n6 vinn.t7 15.0005
R1690 vinn.n22 vinn.t25 15.0005
R1691 vinn.n23 vinn.t6 15.0005
R1692 vinn.n24 vinn.t31 15.0005
R1693 vinn.n25 vinn.t3 15.0005
R1694 vinn.n26 vinn.t30 15.0005
R1695 vinn.n27 vinn.t1 15.0005
R1696 vinn.n28 vinn.t17 15.0005
R1697 vinn vinn.n30 11.8039
R1698 vinn.n29 vinn 10.6252
R1699 vinn.n14 vinn 10.3506
R1700 vinn.n14 vinn 9.95612
R1701 vinn.n29 vinn 9.68456
R1702 vinn vinn.n21 4.90238
R1703 vinn vinn.n13 4.90238
R1704 vinn.n1 vinn.n0 0.6055
R1705 vinn.n2 vinn.n1 0.6055
R1706 vinn.n3 vinn.n2 0.6055
R1707 vinn.n4 vinn.n3 0.6055
R1708 vinn.n5 vinn.n4 0.6055
R1709 vinn.n6 vinn.n5 0.6055
R1710 vinn.n23 vinn.n22 0.6055
R1711 vinn.n24 vinn.n23 0.6055
R1712 vinn.n25 vinn.n24 0.6055
R1713 vinn.n26 vinn.n25 0.6055
R1714 vinn.n27 vinn.n26 0.6055
R1715 vinn.n28 vinn.n27 0.6055
R1716 vinn.n16 vinn.n15 0.6055
R1717 vinn.n17 vinn.n16 0.6055
R1718 vinn.n18 vinn.n17 0.6055
R1719 vinn.n19 vinn.n18 0.6055
R1720 vinn.n20 vinn.n19 0.6055
R1721 vinn.n21 vinn.n20 0.6055
R1722 vinn.n8 vinn.n7 0.6055
R1723 vinn.n9 vinn.n8 0.6055
R1724 vinn.n10 vinn.n9 0.6055
R1725 vinn.n11 vinn.n10 0.6055
R1726 vinn.n12 vinn.n11 0.6055
R1727 vinn.n13 vinn.n12 0.6055
R1728 vinn.n30 vinn.n14 0.548224
R1729 vinn.n30 vinn.n29 0.364638
R1730 vinn vinn.n6 0.333938
R1731 vinn vinn.n28 0.333938
R1732 vout.n15 vout.t12 18.8648
R1733 vout.n7 vout.t16 18.8648
R1734 vout.n11 vout.t13 18.6205
R1735 vout.n4 vout.t9 18.6175
R1736 vout.n17 vout.t19 18.13
R1737 vout.n16 vout.t14 18.13
R1738 vout.n15 vout.t11 18.13
R1739 vout.n9 vout.t10 18.13
R1740 vout.n8 vout.t4 18.13
R1741 vout.n7 vout.t5 18.13
R1742 vout.n13 vout.t15 17.8857
R1743 vout.n12 vout.t17 17.8857
R1744 vout.n11 vout.t6 17.8857
R1745 vout.n6 vout.t7 17.8827
R1746 vout.n5 vout.t8 17.8827
R1747 vout.n4 vout.t18 17.8827
R1748 vout.n3 vout.n2 15.106
R1749 vout.n2 vout.n0 13.7009
R1750 vout.n18 vout.n17 13.4665
R1751 vout.n10 vout.n9 13.4665
R1752 vout.n10 vout.n6 11.8385
R1753 vout.n0 vout.t1 11.1117
R1754 vout.n1 vout.t3 11.1117
R1755 vout.n3 vout 10.8815
R1756 vout.n14 vout.n13 10.3689
R1757 vout.n0 vout.t2 10.2104
R1758 vout.n1 vout.t0 10.2104
R1759 vout.n2 vout.n1 9.36767
R1760 vout.n18 vout.n14 1.4591
R1761 vout vout.n3 0.8673
R1762 vout.n14 vout.n10 0.7507
R1763 vout.n16 vout.n15 0.7353
R1764 vout.n17 vout.n16 0.7353
R1765 vout.n12 vout.n11 0.7353
R1766 vout.n13 vout.n12 0.7353
R1767 vout.n8 vout.n7 0.7353
R1768 vout.n9 vout.n8 0.7353
R1769 vout.n5 vout.n4 0.7353
R1770 vout.n6 vout.n5 0.7353
R1771 vout vout.n18 0.3041
R1772 vdda.n459 vdda.n12 17.0005
R1773 vdda.n459 vdda.n32 17.0005
R1774 vdda.n460 vdda.n459 17.0005
R1775 vdda.n459 vdda.n38 17.0005
R1776 vdda.n459 vdda.n34 17.0005
R1777 vdda.n459 vdda.n35 17.0005
R1778 vdda.n317 vdda.n316 17.0005
R1779 vdda.n318 vdda.n317 17.0005
R1780 vdda.n332 vdda.n331 17.0005
R1781 vdda.n333 vdda.n332 17.0005
R1782 vdda.n347 vdda.n346 17.0005
R1783 vdda.n348 vdda.n347 17.0005
R1784 vdda.n362 vdda.n361 17.0005
R1785 vdda.n363 vdda.n362 17.0005
R1786 vdda.n377 vdda.n376 17.0005
R1787 vdda.n376 vdda.n305 17.0005
R1788 vdda.n384 vdda.n303 17.0005
R1789 vdda.n384 vdda.n383 17.0005
R1790 vdda.n454 vdda.n453 17.0005
R1791 vdda.n453 vdda.n100 17.0005
R1792 vdda.n300 vdda.n195 17.0005
R1793 vdda.n300 vdda.n299 17.0005
R1794 vdda.n291 vdda.n290 17.0005
R1795 vdda.n290 vdda.n289 17.0005
R1796 vdda.n281 vdda.n280 17.0005
R1797 vdda.n280 vdda.n279 17.0005
R1798 vdda.n271 vdda.n270 17.0005
R1799 vdda.n270 vdda.n269 17.0005
R1800 vdda.n261 vdda.n260 17.0005
R1801 vdda.n260 vdda.n259 17.0005
R1802 vdda.n257 vdda.n5 17.0005
R1803 vdda.n6 vdda.n5 17.0005
R1804 vdda.t0 vdda.n104 8.501
R1805 vdda.t0 vdda.n107 8.501
R1806 vdda.t0 vdda.n110 8.501
R1807 vdda.t0 vdda.n113 8.501
R1808 vdda.t0 vdda.n117 8.501
R1809 vdda.t0 vdda.n120 8.501
R1810 vdda.t0 vdda.n123 8.501
R1811 vdda.t0 vdda.n126 8.501
R1812 vdda.t0 vdda.n129 8.501
R1813 vdda.t0 vdda.n132 8.501
R1814 vdda.t0 vdda.n135 8.501
R1815 vdda.t0 vdda.n138 8.501
R1816 vdda.t0 vdda.n141 8.501
R1817 vdda.t0 vdda.n144 8.501
R1818 vdda.t0 vdda.n147 8.501
R1819 vdda.t0 vdda.n150 8.501
R1820 vdda.t0 vdda.n153 8.501
R1821 vdda.t0 vdda.n156 8.501
R1822 vdda.t0 vdda.n159 8.501
R1823 vdda.t0 vdda.n162 8.501
R1824 vdda.t0 vdda.n165 8.501
R1825 vdda.t0 vdda.n168 8.501
R1826 vdda.t0 vdda.n171 8.501
R1827 vdda.t0 vdda.n174 8.501
R1828 vdda.t0 vdda.n177 8.501
R1829 vdda.t0 vdda.n180 8.501
R1830 vdda.t0 vdda.n183 8.501
R1831 vdda.t0 vdda.n186 8.501
R1832 vdda.t0 vdda.n189 8.501
R1833 vdda.t0 vdda.n192 8.501
R1834 vdda.t0 vdda.n385 8.501
R1835 vdda.t0 vdda.n388 8.501
R1836 vdda.t0 vdda.n389 8.501
R1837 vdda.t0 vdda.n93 8.501
R1838 vdda.n452 vdda.t0 8.501
R1839 vdda.t0 vdda.n301 8.501
R1840 vdda.t0 vdda.n191 8.501
R1841 vdda.t0 vdda.n188 8.501
R1842 vdda.t0 vdda.n185 8.501
R1843 vdda.t0 vdda.n182 8.501
R1844 vdda.t0 vdda.n179 8.501
R1845 vdda.t0 vdda.n176 8.501
R1846 vdda.t0 vdda.n173 8.501
R1847 vdda.t0 vdda.n170 8.501
R1848 vdda.t0 vdda.n167 8.501
R1849 vdda.t0 vdda.n164 8.501
R1850 vdda.t0 vdda.n161 8.501
R1851 vdda.t0 vdda.n158 8.501
R1852 vdda.t0 vdda.n155 8.501
R1853 vdda.t0 vdda.n152 8.501
R1854 vdda.t0 vdda.n149 8.501
R1855 vdda.t0 vdda.n146 8.501
R1856 vdda.t0 vdda.n143 8.501
R1857 vdda.t0 vdda.n140 8.501
R1858 vdda.t0 vdda.n137 8.501
R1859 vdda.t0 vdda.n134 8.501
R1860 vdda.t0 vdda.n131 8.501
R1861 vdda.t0 vdda.n128 8.501
R1862 vdda.t0 vdda.n125 8.501
R1863 vdda.t0 vdda.n122 8.501
R1864 vdda.t0 vdda.n119 8.501
R1865 vdda.t0 vdda.n116 8.501
R1866 vdda.t0 vdda.n112 8.501
R1867 vdda.t0 vdda.n109 8.501
R1868 vdda.t0 vdda.n106 8.501
R1869 vdda.t0 vdda.n103 8.501
R1870 vdda.t0 vdda.n451 8.501
R1871 vdda.t0 vdda.n386 8.501
R1872 vdda.t0 vdda.n193 8.501
R1873 vdda.t0 vdda.n190 8.501
R1874 vdda.t0 vdda.n187 8.501
R1875 vdda.t0 vdda.n184 8.501
R1876 vdda.t0 vdda.n181 8.501
R1877 vdda.t0 vdda.n178 8.501
R1878 vdda.t0 vdda.n175 8.501
R1879 vdda.t0 vdda.n172 8.501
R1880 vdda.t0 vdda.n169 8.501
R1881 vdda.t0 vdda.n166 8.501
R1882 vdda.t0 vdda.n163 8.501
R1883 vdda.t0 vdda.n160 8.501
R1884 vdda.t0 vdda.n157 8.501
R1885 vdda.t0 vdda.n154 8.501
R1886 vdda.t0 vdda.n151 8.501
R1887 vdda.t0 vdda.n148 8.501
R1888 vdda.t0 vdda.n145 8.501
R1889 vdda.t0 vdda.n142 8.501
R1890 vdda.t0 vdda.n139 8.501
R1891 vdda.t0 vdda.n136 8.501
R1892 vdda.t0 vdda.n133 8.501
R1893 vdda.t0 vdda.n130 8.501
R1894 vdda.t0 vdda.n127 8.501
R1895 vdda.t0 vdda.n124 8.501
R1896 vdda.t0 vdda.n121 8.501
R1897 vdda.t0 vdda.n118 8.501
R1898 vdda.t0 vdda.n115 8.501
R1899 vdda.t0 vdda.n111 8.501
R1900 vdda.t0 vdda.n108 8.501
R1901 vdda.t0 vdda.n105 8.501
R1902 vdda.t0 vdda.n102 8.501
R1903 vdda.n315 vdda.n314 8.46995
R1904 vdda.n320 vdda.n319 8.46995
R1905 vdda.n322 vdda.n321 8.46995
R1906 vdda.n324 vdda.n323 8.46995
R1907 vdda.n326 vdda.n325 8.46995
R1908 vdda.n328 vdda.n327 8.46995
R1909 vdda.n330 vdda.n329 8.46995
R1910 vdda.n335 vdda.n334 8.46995
R1911 vdda.n337 vdda.n336 8.46995
R1912 vdda.n339 vdda.n338 8.46995
R1913 vdda.n341 vdda.n340 8.46995
R1914 vdda.n343 vdda.n342 8.46995
R1915 vdda.n345 vdda.n344 8.46995
R1916 vdda.n350 vdda.n349 8.46995
R1917 vdda.n352 vdda.n351 8.46995
R1918 vdda.n354 vdda.n353 8.46995
R1919 vdda.n356 vdda.n355 8.46995
R1920 vdda.n358 vdda.n357 8.46995
R1921 vdda.n360 vdda.n359 8.46995
R1922 vdda.n365 vdda.n364 8.46995
R1923 vdda.n367 vdda.n366 8.46995
R1924 vdda.n369 vdda.n368 8.46995
R1925 vdda.n371 vdda.n370 8.46995
R1926 vdda.n373 vdda.n372 8.46995
R1927 vdda.n375 vdda.n374 8.46995
R1928 vdda.n304 vdda.n302 8.46995
R1929 vdda.n392 vdda.n391 8.46995
R1930 vdda.n393 vdda.n390 8.46995
R1931 vdda.n459 vdda.n458 8.46995
R1932 vdda.n457 vdda.n95 8.46995
R1933 vdda.n194 vdda.n101 8.46995
R1934 vdda.n298 vdda.n197 8.46995
R1935 vdda.n297 vdda.n198 8.46995
R1936 vdda.n296 vdda.n199 8.46995
R1937 vdda.n294 vdda.n201 8.46995
R1938 vdda.n293 vdda.n202 8.46995
R1939 vdda.n292 vdda.n203 8.46995
R1940 vdda.n288 vdda.n205 8.46995
R1941 vdda.n287 vdda.n206 8.46995
R1942 vdda.n286 vdda.n207 8.46995
R1943 vdda.n284 vdda.n209 8.46995
R1944 vdda.n283 vdda.n210 8.46995
R1945 vdda.n282 vdda.n211 8.46995
R1946 vdda.n278 vdda.n213 8.46995
R1947 vdda.n277 vdda.n214 8.46995
R1948 vdda.n276 vdda.n215 8.46995
R1949 vdda.n274 vdda.n217 8.46995
R1950 vdda.n273 vdda.n218 8.46995
R1951 vdda.n272 vdda.n219 8.46995
R1952 vdda.n268 vdda.n221 8.46995
R1953 vdda.n267 vdda.n222 8.46995
R1954 vdda.n266 vdda.n223 8.46995
R1955 vdda.n264 vdda.n225 8.46995
R1956 vdda.n263 vdda.n226 8.46995
R1957 vdda.n262 vdda.n227 8.46995
R1958 vdda.n258 vdda.n229 8.46995
R1959 vdda.n447 vdda.n394 8.46995
R1960 vdda.n446 vdda.n395 8.46995
R1961 vdda.n445 vdda.n396 8.46995
R1962 vdda.n444 vdda.n397 8.46995
R1963 vdda.n443 vdda.n398 8.46995
R1964 vdda.n442 vdda.n399 8.46995
R1965 vdda.n441 vdda.n400 8.46995
R1966 vdda.n440 vdda.n401 8.46995
R1967 vdda.n439 vdda.n402 8.46995
R1968 vdda.n438 vdda.n403 8.46995
R1969 vdda.n437 vdda.n404 8.46995
R1970 vdda.n436 vdda.n405 8.46995
R1971 vdda.n435 vdda.n406 8.46995
R1972 vdda.n434 vdda.n407 8.46995
R1973 vdda.n433 vdda.n408 8.46995
R1974 vdda.n432 vdda.n409 8.46995
R1975 vdda.n431 vdda.n410 8.46995
R1976 vdda.n430 vdda.n411 8.46995
R1977 vdda.n429 vdda.n412 8.46995
R1978 vdda.n428 vdda.n413 8.46995
R1979 vdda.n427 vdda.n414 8.46995
R1980 vdda.n426 vdda.n415 8.46995
R1981 vdda.n425 vdda.n416 8.46995
R1982 vdda.n424 vdda.n417 8.46995
R1983 vdda.n423 vdda.n418 8.46995
R1984 vdda.n422 vdda.n419 8.46995
R1985 vdda.n421 vdda.n420 8.46995
R1986 vdda.n114 vdda.n0 8.46995
R1987 vdda.n467 vdda.n1 8.46995
R1988 vdda.n466 vdda.n2 8.46995
R1989 vdda.n465 vdda.n3 8.46995
R1990 vdda.n464 vdda.n4 8.46995
R1991 vdda.n87 vdda.t36 7.44301
R1992 vdda.n69 vdda.t66 7.44301
R1993 vdda.n16 vdda.t19 7.44301
R1994 vdda.n29 vdda.t40 7.44301
R1995 vdda.n311 vdda.t63 7.44301
R1996 vdda.n380 vdda.t34 7.44301
R1997 vdda.n236 vdda.t26 7.44301
R1998 vdda.n254 vdda.t54 7.44301
R1999 vdda.n20 vdda.t7 6.20273
R2000 vdda.n22 vdda.t8 6.20273
R2001 vdda.n24 vdda.t5 6.20273
R2002 vdda.n308 vdda.t4 6.20273
R2003 vdda.n307 vdda.t6 6.20273
R2004 vdda.n306 vdda.t3 6.20273
R2005 vdda.t0 vdda.n387 5.66778
R2006 vdda.t0 vdda.n33 5.66767
R2007 vdda.t0 vdda.n450 5.66767
R2008 vdda.n97 vdda.n96 5.63414
R2009 vdda.n456 vdda.n96 5.61281
R2010 vdda.n449 vdda.n448 5.59203
R2011 vdda.n50 vdda.t23 5.56245
R2012 vdda.n52 vdda.t23 5.56245
R2013 vdda.n54 vdda.t23 5.56245
R2014 vdda.n56 vdda.t23 5.56245
R2015 vdda.n58 vdda.t23 5.56245
R2016 vdda.n60 vdda.t23 5.56245
R2017 vdda.n62 vdda.t23 5.56245
R2018 vdda.n64 vdda.t23 5.56245
R2019 vdda.n66 vdda.t23 5.56245
R2020 vdda.n68 vdda.t68 5.56245
R2021 vdda.n88 vdda.t23 5.56245
R2022 vdda.n15 vdda.t21 5.56245
R2023 vdda.n17 vdda.t2 5.56245
R2024 vdda.n28 vdda.t16 5.56245
R2025 vdda.n30 vdda.t16 5.56245
R2026 vdda.n310 vdda.t65 5.56245
R2027 vdda.n312 vdda.t1 5.56245
R2028 vdda.n379 vdda.t13 5.56245
R2029 vdda.n381 vdda.t13 5.56245
R2030 vdda.t18 vdda.n234 5.56245
R2031 vdda.t18 vdda.n200 5.56245
R2032 vdda.t18 vdda.n233 5.56245
R2033 vdda.t18 vdda.n208 5.56245
R2034 vdda.t18 vdda.n232 5.56245
R2035 vdda.t18 vdda.n216 5.56245
R2036 vdda.t18 vdda.n231 5.56245
R2037 vdda.t18 vdda.n224 5.56245
R2038 vdda.t18 vdda.n230 5.56245
R2039 vdda.n255 vdda.t56 5.56245
R2040 vdda.n235 vdda.t18 5.56245
R2041 vdda.t0 vdda.n99 4.251
R2042 vdda.n459 vdda.n26 4.17429
R2043 vdda.n459 vdda.n48 4.17416
R2044 vdda.n459 vdda.n13 4.17295
R2045 vdda.n459 vdda.n39 4.17282
R2046 vdda.n85 vdda.t59 2.82253
R2047 vdda.n83 vdda.t30 2.82253
R2048 vdda.n81 vdda.t52 2.82253
R2049 vdda.n79 vdda.t38 2.82253
R2050 vdda.n77 vdda.t57 2.82253
R2051 vdda.n75 vdda.t32 2.82253
R2052 vdda.n73 vdda.t50 2.82253
R2053 vdda.n71 vdda.t22 2.82253
R2054 vdda.n238 vdda.t48 2.82253
R2055 vdda.n240 vdda.t17 2.82253
R2056 vdda.n242 vdda.t44 2.82253
R2057 vdda.n244 vdda.t28 2.82253
R2058 vdda.n246 vdda.t46 2.82253
R2059 vdda.n248 vdda.t24 2.82253
R2060 vdda.n250 vdda.t42 2.82253
R2061 vdda.n252 vdda.t61 2.82253
R2062 vdda.n469 vdda.n468 2.55416
R2063 vdda.n463 vdda.n5 2.29632
R2064 vdda.n461 vdda.n5 2.29413
R2065 vdda.n459 vdda.n47 2.29267
R2066 vdda.n459 vdda.n46 2.29267
R2067 vdda.n459 vdda.n45 2.29267
R2068 vdda.n459 vdda.n44 2.29267
R2069 vdda.n459 vdda.n43 2.29267
R2070 vdda.n459 vdda.n42 2.29267
R2071 vdda.n459 vdda.n41 2.29267
R2072 vdda.n459 vdda.n40 2.2913
R2073 vdda.n459 vdda.n9 1.72624
R2074 vdda.n459 vdda.n10 1.72331
R2075 vdda.n459 vdda.n90 1.70496
R2076 vdda.n459 vdda.n92 1.52264
R2077 vdda.n37 vdda 1.205
R2078 vdda.n69 vdda.n68 0.987904
R2079 vdda.n16 vdda.n15 0.987904
R2080 vdda.n17 vdda.n16 0.987904
R2081 vdda.n29 vdda.n28 0.987904
R2082 vdda.n311 vdda.n310 0.987904
R2083 vdda.n312 vdda.n311 0.987904
R2084 vdda.n380 vdda.n379 0.987904
R2085 vdda.n255 vdda.n254 0.987904
R2086 vdda.n88 vdda.n87 0.987558
R2087 vdda.n30 vdda.n29 0.987558
R2088 vdda.n381 vdda.n380 0.987558
R2089 vdda.n236 vdda.n235 0.987558
R2090 vdda.n459 vdda.n21 0.968021
R2091 vdda.n459 vdda.n23 0.968021
R2092 vdda.n459 vdda.n25 0.968021
R2093 vdda.n459 vdda.n19 0.966815
R2094 vdda.n20 vdda.n19 0.810176
R2095 vdda.n27 vdda.n25 0.808344
R2096 vdda.n24 vdda.n23 0.808344
R2097 vdda.n22 vdda.n21 0.808344
R2098 vdda.n85 vdda.n84 0.803704
R2099 vdda.n83 vdda.n82 0.803704
R2100 vdda.n81 vdda.n80 0.803704
R2101 vdda.n79 vdda.n78 0.803704
R2102 vdda.n77 vdda.n76 0.803704
R2103 vdda.n75 vdda.n74 0.803704
R2104 vdda.n73 vdda.n72 0.803704
R2105 vdda.n71 vdda.n70 0.803704
R2106 vdda.n239 vdda.n238 0.803704
R2107 vdda.n241 vdda.n240 0.803704
R2108 vdda.n243 vdda.n242 0.803704
R2109 vdda.n245 vdda.n244 0.803704
R2110 vdda.n247 vdda.n246 0.803704
R2111 vdda.n249 vdda.n248 0.803704
R2112 vdda.n251 vdda.n250 0.803704
R2113 vdda.n253 vdda.n252 0.803704
R2114 vdda.n86 vdda.n85 0.802423
R2115 vdda.n84 vdda.n83 0.802423
R2116 vdda.n82 vdda.n81 0.802423
R2117 vdda.n80 vdda.n79 0.802423
R2118 vdda.n78 vdda.n77 0.802423
R2119 vdda.n76 vdda.n75 0.802423
R2120 vdda.n74 vdda.n73 0.802423
R2121 vdda.n72 vdda.n71 0.802423
R2122 vdda.n238 vdda.n237 0.802423
R2123 vdda.n240 vdda.n239 0.802423
R2124 vdda.n242 vdda.n241 0.802423
R2125 vdda.n244 vdda.n243 0.802423
R2126 vdda.n246 vdda.n245 0.802423
R2127 vdda.n248 vdda.n247 0.802423
R2128 vdda.n250 vdda.n249 0.802423
R2129 vdda.n252 vdda.n251 0.802423
R2130 vdda.n25 vdda.n24 0.767309
R2131 vdda.n23 vdda.n22 0.767309
R2132 vdda.n21 vdda.n20 0.767309
R2133 vdda.n19 vdda.n18 0.763505
R2134 vdda.n50 vdda.n49 0.64112
R2135 vdda.n52 vdda.n51 0.64112
R2136 vdda.n54 vdda.n53 0.64112
R2137 vdda.n56 vdda.n55 0.64112
R2138 vdda.n58 vdda.n57 0.64112
R2139 vdda.n60 vdda.n59 0.64112
R2140 vdda.n62 vdda.n61 0.64112
R2141 vdda.n64 vdda.n63 0.64112
R2142 vdda.n89 vdda.n88 0.64112
R2143 vdda.n31 vdda.n30 0.64112
R2144 vdda.n382 vdda.n381 0.64112
R2145 vdda.n234 vdda.n196 0.64112
R2146 vdda.n295 vdda.n200 0.64112
R2147 vdda.n233 vdda.n204 0.64112
R2148 vdda.n285 vdda.n208 0.64112
R2149 vdda.n232 vdda.n212 0.64112
R2150 vdda.n275 vdda.n216 0.64112
R2151 vdda.n231 vdda.n220 0.64112
R2152 vdda.n265 vdda.n224 0.64112
R2153 vdda.n235 vdda.n98 0.64112
R2154 vdda.n66 vdda.n65 0.640774
R2155 vdda.n68 vdda.n67 0.640774
R2156 vdda.n15 vdda.n14 0.640774
R2157 vdda.n18 vdda.n17 0.640774
R2158 vdda.n28 vdda.n27 0.640774
R2159 vdda.n310 vdda.n309 0.640774
R2160 vdda.n313 vdda.n312 0.640774
R2161 vdda.n379 vdda.n378 0.640774
R2162 vdda.n230 vdda.n228 0.640774
R2163 vdda.n256 vdda.n255 0.640774
R2164 vdda.n90 vdda.n89 0.636597
R2165 vdda.n11 vdda.n9 0.552389
R2166 vdda.n91 vdda.n90 0.543067
R2167 vdda.n37 vdda.n10 0.522655
R2168 vdda.n70 vdda.n66 0.513933
R2169 vdda.n253 vdda.n230 0.513933
R2170 vdda.n86 vdda.n50 0.513587
R2171 vdda.n84 vdda.n52 0.513587
R2172 vdda.n82 vdda.n54 0.513587
R2173 vdda.n80 vdda.n56 0.513587
R2174 vdda.n78 vdda.n58 0.513587
R2175 vdda.n76 vdda.n60 0.513587
R2176 vdda.n74 vdda.n62 0.513587
R2177 vdda.n72 vdda.n64 0.513587
R2178 vdda.n237 vdda.n234 0.513587
R2179 vdda.n239 vdda.n200 0.513587
R2180 vdda.n241 vdda.n233 0.513587
R2181 vdda.n243 vdda.n208 0.513587
R2182 vdda.n245 vdda.n232 0.513587
R2183 vdda.n247 vdda.n216 0.513587
R2184 vdda.n249 vdda.n231 0.513587
R2185 vdda.n251 vdda.n224 0.513587
R2186 vdda.n92 vdda.n91 0.487895
R2187 vdda.n461 vdda.n460 0.487765
R2188 vdda.n87 vdda.n86 0.474471
R2189 vdda.n70 vdda.n69 0.474471
R2190 vdda.n237 vdda.n236 0.474471
R2191 vdda.n254 vdda.n253 0.474471
R2192 vdda.n63 vdda.n40 0.454505
R2193 vdda.n49 vdda.n47 0.4496
R2194 vdda.n51 vdda.n46 0.4496
R2195 vdda.n53 vdda.n45 0.4496
R2196 vdda.n55 vdda.n44 0.4496
R2197 vdda.n57 vdda.n43 0.4496
R2198 vdda.n59 vdda.n42 0.4496
R2199 vdda.n61 vdda.n41 0.4496
R2200 vdda.n94 vdda.n92 0.438254
R2201 vdda.n11 vdda.n10 0.416748
R2202 vdda.n51 vdda.n47 0.405126
R2203 vdda.n53 vdda.n46 0.405126
R2204 vdda.n55 vdda.n45 0.405126
R2205 vdda.n57 vdda.n44 0.405126
R2206 vdda.n59 vdda.n43 0.405126
R2207 vdda.n61 vdda.n42 0.405126
R2208 vdda.n63 vdda.n41 0.405126
R2209 vdda.n65 vdda.n40 0.399705
R2210 vdda.n9 vdda.n7 0.388549
R2211 vdda.n463 vdda.n462 0.388318
R2212 vdda vdda.n463 0.381578
R2213 vdda.n462 vdda.n461 0.354662
R2214 vdda.n448 vdda.n447 0.343481
R2215 vdda.n448 vdda.n393 0.342175
R2216 vdda.n457 vdda.n456 0.312698
R2217 vdda.n65 vdda.n39 0.283787
R2218 vdda.n18 vdda.n13 0.283654
R2219 vdda.n392 vdda.n97 0.280735
R2220 vdda.n89 vdda.n48 0.278395
R2221 vdda.n31 vdda.n26 0.278262
R2222 vdda.n324 vdda.n322 0.257711
R2223 vdda.n264 vdda.n263 0.257711
R2224 vdda.n421 vdda.n0 0.257711
R2225 vdda.n466 vdda.n465 0.257711
R2226 vdda.n375 vdda.n373 0.250378
R2227 vdda.n373 vdda.n371 0.250378
R2228 vdda.n371 vdda.n369 0.250378
R2229 vdda.n369 vdda.n367 0.250378
R2230 vdda.n367 vdda.n365 0.250378
R2231 vdda.n360 vdda.n358 0.250378
R2232 vdda.n358 vdda.n356 0.250378
R2233 vdda.n356 vdda.n354 0.250378
R2234 vdda.n354 vdda.n352 0.250378
R2235 vdda.n352 vdda.n350 0.250378
R2236 vdda.n345 vdda.n343 0.250378
R2237 vdda.n343 vdda.n341 0.250378
R2238 vdda.n341 vdda.n339 0.250378
R2239 vdda.n339 vdda.n337 0.250378
R2240 vdda.n337 vdda.n335 0.250378
R2241 vdda.n330 vdda.n328 0.250378
R2242 vdda.n328 vdda.n326 0.250378
R2243 vdda.n326 vdda.n324 0.250378
R2244 vdda.n322 vdda.n320 0.250378
R2245 vdda.n393 vdda.n392 0.250378
R2246 vdda.n458 vdda.n457 0.250378
R2247 vdda.n298 vdda.n297 0.250378
R2248 vdda.n297 vdda.n296 0.250378
R2249 vdda.n294 vdda.n293 0.250378
R2250 vdda.n293 vdda.n292 0.250378
R2251 vdda.n288 vdda.n287 0.250378
R2252 vdda.n287 vdda.n286 0.250378
R2253 vdda.n284 vdda.n283 0.250378
R2254 vdda.n283 vdda.n282 0.250378
R2255 vdda.n278 vdda.n277 0.250378
R2256 vdda.n277 vdda.n276 0.250378
R2257 vdda.n274 vdda.n273 0.250378
R2258 vdda.n273 vdda.n272 0.250378
R2259 vdda.n268 vdda.n267 0.250378
R2260 vdda.n267 vdda.n266 0.250378
R2261 vdda.n263 vdda.n262 0.250378
R2262 vdda.n447 vdda.n446 0.250378
R2263 vdda.n446 vdda.n445 0.250378
R2264 vdda.n445 vdda.n444 0.250378
R2265 vdda.n444 vdda.n443 0.250378
R2266 vdda.n443 vdda.n442 0.250378
R2267 vdda.n442 vdda.n441 0.250378
R2268 vdda.n441 vdda.n440 0.250378
R2269 vdda.n440 vdda.n439 0.250378
R2270 vdda.n439 vdda.n438 0.250378
R2271 vdda.n438 vdda.n437 0.250378
R2272 vdda.n437 vdda.n436 0.250378
R2273 vdda.n436 vdda.n435 0.250378
R2274 vdda.n435 vdda.n434 0.250378
R2275 vdda.n434 vdda.n433 0.250378
R2276 vdda.n433 vdda.n432 0.250378
R2277 vdda.n432 vdda.n431 0.250378
R2278 vdda.n431 vdda.n430 0.250378
R2279 vdda.n430 vdda.n429 0.250378
R2280 vdda.n429 vdda.n428 0.250378
R2281 vdda.n428 vdda.n427 0.250378
R2282 vdda.n427 vdda.n426 0.250378
R2283 vdda.n426 vdda.n425 0.250378
R2284 vdda.n425 vdda.n424 0.250378
R2285 vdda.n424 vdda.n423 0.250378
R2286 vdda.n423 vdda.n422 0.250378
R2287 vdda.n422 vdda.n421 0.250378
R2288 vdda.n467 vdda.n466 0.250378
R2289 vdda.n465 vdda.n464 0.250378
R2290 vdda.n456 vdda.n455 0.236919
R2291 vdda.n27 vdda.n26 0.227191
R2292 vdda.n49 vdda.n48 0.227062
R2293 vdda.n14 vdda.n13 0.221637
R2294 vdda.n67 vdda.n39 0.221508
R2295 vdda.n91 vdda.n32 0.2205
R2296 vdda.n383 vdda.n94 0.2205
R2297 vdda.n455 vdda.n454 0.2205
R2298 vdda.t0 vdda.n36 0.201
R2299 vdda.n316 vdda.n315 0.195106
R2300 vdda.n259 vdda.n258 0.195106
R2301 vdda.n304 vdda.n303 0.187772
R2302 vdda.n305 vdda.n304 0.187772
R2303 vdda.n377 vdda.n375 0.187772
R2304 vdda.n365 vdda.n363 0.187772
R2305 vdda.n361 vdda.n360 0.187772
R2306 vdda.n350 vdda.n348 0.187772
R2307 vdda.n346 vdda.n345 0.187772
R2308 vdda.n335 vdda.n333 0.187772
R2309 vdda.n331 vdda.n330 0.187772
R2310 vdda.n320 vdda.n318 0.187772
R2311 vdda.n315 vdda.n35 0.187772
R2312 vdda.n194 vdda.n100 0.187772
R2313 vdda.n195 vdda.n194 0.187772
R2314 vdda.n299 vdda.n298 0.187772
R2315 vdda.n292 vdda.n291 0.187772
R2316 vdda.n289 vdda.n288 0.187772
R2317 vdda.n282 vdda.n281 0.187772
R2318 vdda.n279 vdda.n278 0.187772
R2319 vdda.n272 vdda.n271 0.187772
R2320 vdda.n269 vdda.n268 0.187772
R2321 vdda.n262 vdda.n261 0.187772
R2322 vdda.n258 vdda.n257 0.187772
R2323 vdda.n458 vdda.n94 0.182272
R2324 vdda.n464 vdda 0.180439
R2325 vdda.t0 vdda.n8 0.171785
R2326 vdda.n38 vdda.n37 0.161833
R2327 vdda.n12 vdda.n11 0.161833
R2328 vdda.n34 vdda.n7 0.161833
R2329 vdda.n462 vdda.n6 0.161833
R2330 vdda.n468 vdda.n0 0.160272
R2331 vdda.n295 vdda.n294 0.147439
R2332 vdda.n285 vdda.n284 0.147439
R2333 vdda.n275 vdda.n274 0.147439
R2334 vdda.n265 vdda.n264 0.147439
R2335 vdda.n460 vdda.n7 0.119667
R2336 vdda.n296 vdda.n295 0.103439
R2337 vdda.n286 vdda.n285 0.103439
R2338 vdda.n276 vdda.n275 0.103439
R2339 vdda.n266 vdda.n265 0.103439
R2340 vdda.n67 vdda.n38 0.0921667
R2341 vdda.n14 vdda.n12 0.0921667
R2342 vdda.n382 vdda.n303 0.0921667
R2343 vdda.n316 vdda.n313 0.0921667
R2344 vdda.n309 vdda.n34 0.0921667
R2345 vdda.n100 vdda.n98 0.0921667
R2346 vdda.n259 vdda.n228 0.0921667
R2347 vdda.n256 vdda.n6 0.0921667
R2348 vdda.n468 vdda.n467 0.0906056
R2349 vdda.n378 vdda.n377 0.0848333
R2350 vdda.n361 vdda.n306 0.0848333
R2351 vdda.n346 vdda.n307 0.0848333
R2352 vdda.n331 vdda.n308 0.0848333
R2353 vdda.n299 vdda.n196 0.0848333
R2354 vdda.n289 vdda.n204 0.0848333
R2355 vdda.n279 vdda.n212 0.0848333
R2356 vdda.n269 vdda.n220 0.0848333
R2357 vdda.n455 vdda.n97 0.0609304
R2358 vdda.n378 vdda.n305 0.0408333
R2359 vdda.n363 vdda.n306 0.0408333
R2360 vdda.n348 vdda.n307 0.0408333
R2361 vdda.n333 vdda.n308 0.0408333
R2362 vdda.n196 vdda.n195 0.0408333
R2363 vdda.n291 vdda.n204 0.0408333
R2364 vdda.n281 vdda.n212 0.0408333
R2365 vdda.n271 vdda.n220 0.0408333
R2366 vdda.n32 vdda.n31 0.0335
R2367 vdda.n383 vdda.n382 0.0335
R2368 vdda.n318 vdda.n313 0.0335
R2369 vdda.n309 vdda.n35 0.0335
R2370 vdda.n454 vdda.n98 0.0335
R2371 vdda.n261 vdda.n228 0.0335
R2372 vdda.n257 vdda.n256 0.0335
R2373 vdda.n469 vdda 0.0151933
R2374 vdda vdda.n469 0.0140551
R2375 vdda.n459 vdda.n8 0.0020653
R2376 vdda.n8 vdda.n5 0.0019343
R2377 vdda.n387 vdda.n95 0.00166667
R2378 vdda.n387 vdda.n96 0.00133332
R2379 vdda.n459 vdda.n36 0.001
R2380 vdda.n384 vdda.n36 0.001
R2381 vdda.n385 vdda.n302 0.001
R2382 vdda.n376 vdda.n192 0.001
R2383 vdda.n374 vdda.n189 0.001
R2384 vdda.n372 vdda.n186 0.001
R2385 vdda.n370 vdda.n183 0.001
R2386 vdda.n368 vdda.n180 0.001
R2387 vdda.n366 vdda.n177 0.001
R2388 vdda.n364 vdda.n174 0.001
R2389 vdda.n362 vdda.n171 0.001
R2390 vdda.n359 vdda.n168 0.001
R2391 vdda.n357 vdda.n165 0.001
R2392 vdda.n355 vdda.n162 0.001
R2393 vdda.n353 vdda.n159 0.001
R2394 vdda.n351 vdda.n156 0.001
R2395 vdda.n349 vdda.n153 0.001
R2396 vdda.n347 vdda.n150 0.001
R2397 vdda.n344 vdda.n147 0.001
R2398 vdda.n342 vdda.n144 0.001
R2399 vdda.n340 vdda.n141 0.001
R2400 vdda.n338 vdda.n138 0.001
R2401 vdda.n336 vdda.n135 0.001
R2402 vdda.n334 vdda.n132 0.001
R2403 vdda.n332 vdda.n129 0.001
R2404 vdda.n329 vdda.n126 0.001
R2405 vdda.n327 vdda.n123 0.001
R2406 vdda.n325 vdda.n120 0.001
R2407 vdda.n323 vdda.n117 0.001
R2408 vdda.n321 vdda.n113 0.001
R2409 vdda.n319 vdda.n110 0.001
R2410 vdda.n317 vdda.n107 0.001
R2411 vdda.n314 vdda.n104 0.001
R2412 vdda.n314 vdda.n33 0.001
R2413 vdda.n459 vdda.n33 0.001
R2414 vdda.n317 vdda.n104 0.001
R2415 vdda.n319 vdda.n107 0.001
R2416 vdda.n321 vdda.n110 0.001
R2417 vdda.n323 vdda.n113 0.001
R2418 vdda.n325 vdda.n117 0.001
R2419 vdda.n327 vdda.n120 0.001
R2420 vdda.n329 vdda.n123 0.001
R2421 vdda.n332 vdda.n126 0.001
R2422 vdda.n334 vdda.n129 0.001
R2423 vdda.n336 vdda.n132 0.001
R2424 vdda.n338 vdda.n135 0.001
R2425 vdda.n340 vdda.n138 0.001
R2426 vdda.n342 vdda.n141 0.001
R2427 vdda.n344 vdda.n144 0.001
R2428 vdda.n347 vdda.n147 0.001
R2429 vdda.n349 vdda.n150 0.001
R2430 vdda.n351 vdda.n153 0.001
R2431 vdda.n353 vdda.n156 0.001
R2432 vdda.n355 vdda.n159 0.001
R2433 vdda.n357 vdda.n162 0.001
R2434 vdda.n359 vdda.n165 0.001
R2435 vdda.n362 vdda.n168 0.001
R2436 vdda.n364 vdda.n171 0.001
R2437 vdda.n366 vdda.n174 0.001
R2438 vdda.n368 vdda.n177 0.001
R2439 vdda.n370 vdda.n180 0.001
R2440 vdda.n372 vdda.n183 0.001
R2441 vdda.n374 vdda.n186 0.001
R2442 vdda.n376 vdda.n189 0.001
R2443 vdda.n302 vdda.n192 0.001
R2444 vdda.n385 vdda.n384 0.001
R2445 vdda.n459 vdda.n93 0.001
R2446 vdda.n453 vdda.n99 0.001
R2447 vdda.n452 vdda.n101 0.001
R2448 vdda.n301 vdda.n300 0.001
R2449 vdda.n197 vdda.n191 0.001
R2450 vdda.n198 vdda.n188 0.001
R2451 vdda.n199 vdda.n185 0.001
R2452 vdda.n201 vdda.n182 0.001
R2453 vdda.n202 vdda.n179 0.001
R2454 vdda.n203 vdda.n176 0.001
R2455 vdda.n290 vdda.n173 0.001
R2456 vdda.n205 vdda.n170 0.001
R2457 vdda.n206 vdda.n167 0.001
R2458 vdda.n207 vdda.n164 0.001
R2459 vdda.n209 vdda.n161 0.001
R2460 vdda.n210 vdda.n158 0.001
R2461 vdda.n211 vdda.n155 0.001
R2462 vdda.n280 vdda.n152 0.001
R2463 vdda.n213 vdda.n149 0.001
R2464 vdda.n214 vdda.n146 0.001
R2465 vdda.n215 vdda.n143 0.001
R2466 vdda.n217 vdda.n140 0.001
R2467 vdda.n218 vdda.n137 0.001
R2468 vdda.n219 vdda.n134 0.001
R2469 vdda.n270 vdda.n131 0.001
R2470 vdda.n221 vdda.n128 0.001
R2471 vdda.n222 vdda.n125 0.001
R2472 vdda.n223 vdda.n122 0.001
R2473 vdda.n225 vdda.n119 0.001
R2474 vdda.n226 vdda.n116 0.001
R2475 vdda.n227 vdda.n112 0.001
R2476 vdda.n260 vdda.n109 0.001
R2477 vdda.n229 vdda.n106 0.001
R2478 vdda.n103 vdda.n5 0.001
R2479 vdda.n394 vdda.n386 0.001
R2480 vdda.n395 vdda.n193 0.001
R2481 vdda.n396 vdda.n190 0.001
R2482 vdda.n397 vdda.n187 0.001
R2483 vdda.n398 vdda.n184 0.001
R2484 vdda.n399 vdda.n181 0.001
R2485 vdda.n400 vdda.n178 0.001
R2486 vdda.n401 vdda.n175 0.001
R2487 vdda.n402 vdda.n172 0.001
R2488 vdda.n403 vdda.n169 0.001
R2489 vdda.n404 vdda.n166 0.001
R2490 vdda.n405 vdda.n163 0.001
R2491 vdda.n406 vdda.n160 0.001
R2492 vdda.n407 vdda.n157 0.001
R2493 vdda.n408 vdda.n154 0.001
R2494 vdda.n409 vdda.n151 0.001
R2495 vdda.n410 vdda.n148 0.001
R2496 vdda.n411 vdda.n145 0.001
R2497 vdda.n412 vdda.n142 0.001
R2498 vdda.n413 vdda.n139 0.001
R2499 vdda.n414 vdda.n136 0.001
R2500 vdda.n415 vdda.n133 0.001
R2501 vdda.n416 vdda.n130 0.001
R2502 vdda.n417 vdda.n127 0.001
R2503 vdda.n418 vdda.n124 0.001
R2504 vdda.n419 vdda.n121 0.001
R2505 vdda.n420 vdda.n118 0.001
R2506 vdda.n115 vdda.n114 0.001
R2507 vdda.n111 vdda.n1 0.001
R2508 vdda.n108 vdda.n2 0.001
R2509 vdda.n105 vdda.n3 0.001
R2510 vdda.n102 vdda.n4 0.001
R2511 vdda.n451 vdda.n5 0.001
R2512 vdda.n388 vdda.n96 0.001
R2513 vdda.n391 vdda.n389 0.001
R2514 vdda.n450 vdda.n390 0.001
R2515 vdda.n391 vdda.n388 0.001
R2516 vdda.n390 vdda.n389 0.001
R2517 vdda.n95 vdda.n93 0.001
R2518 vdda.n99 vdda.n96 0.001
R2519 vdda.n453 vdda.n452 0.001
R2520 vdda.n301 vdda.n101 0.001
R2521 vdda.n300 vdda.n191 0.001
R2522 vdda.n197 vdda.n188 0.001
R2523 vdda.n198 vdda.n185 0.001
R2524 vdda.n199 vdda.n182 0.001
R2525 vdda.n201 vdda.n179 0.001
R2526 vdda.n202 vdda.n176 0.001
R2527 vdda.n203 vdda.n173 0.001
R2528 vdda.n290 vdda.n170 0.001
R2529 vdda.n205 vdda.n167 0.001
R2530 vdda.n206 vdda.n164 0.001
R2531 vdda.n207 vdda.n161 0.001
R2532 vdda.n209 vdda.n158 0.001
R2533 vdda.n210 vdda.n155 0.001
R2534 vdda.n211 vdda.n152 0.001
R2535 vdda.n280 vdda.n149 0.001
R2536 vdda.n213 vdda.n146 0.001
R2537 vdda.n214 vdda.n143 0.001
R2538 vdda.n215 vdda.n140 0.001
R2539 vdda.n217 vdda.n137 0.001
R2540 vdda.n218 vdda.n134 0.001
R2541 vdda.n219 vdda.n131 0.001
R2542 vdda.n270 vdda.n128 0.001
R2543 vdda.n221 vdda.n125 0.001
R2544 vdda.n222 vdda.n122 0.001
R2545 vdda.n223 vdda.n119 0.001
R2546 vdda.n225 vdda.n116 0.001
R2547 vdda.n226 vdda.n112 0.001
R2548 vdda.n227 vdda.n109 0.001
R2549 vdda.n260 vdda.n106 0.001
R2550 vdda.n229 vdda.n103 0.001
R2551 vdda.n450 vdda.n449 0.001
R2552 vdda.n449 vdda.n386 0.001
R2553 vdda.n394 vdda.n193 0.001
R2554 vdda.n395 vdda.n190 0.001
R2555 vdda.n396 vdda.n187 0.001
R2556 vdda.n397 vdda.n184 0.001
R2557 vdda.n398 vdda.n181 0.001
R2558 vdda.n399 vdda.n178 0.001
R2559 vdda.n400 vdda.n175 0.001
R2560 vdda.n401 vdda.n172 0.001
R2561 vdda.n402 vdda.n169 0.001
R2562 vdda.n403 vdda.n166 0.001
R2563 vdda.n404 vdda.n163 0.001
R2564 vdda.n405 vdda.n160 0.001
R2565 vdda.n406 vdda.n157 0.001
R2566 vdda.n407 vdda.n154 0.001
R2567 vdda.n408 vdda.n151 0.001
R2568 vdda.n409 vdda.n148 0.001
R2569 vdda.n410 vdda.n145 0.001
R2570 vdda.n411 vdda.n142 0.001
R2571 vdda.n412 vdda.n139 0.001
R2572 vdda.n413 vdda.n136 0.001
R2573 vdda.n414 vdda.n133 0.001
R2574 vdda.n415 vdda.n130 0.001
R2575 vdda.n416 vdda.n127 0.001
R2576 vdda.n417 vdda.n124 0.001
R2577 vdda.n418 vdda.n121 0.001
R2578 vdda.n419 vdda.n118 0.001
R2579 vdda.n420 vdda.n115 0.001
R2580 vdda.n114 vdda.n111 0.001
R2581 vdda.n108 vdda.n1 0.001
R2582 vdda.n105 vdda.n2 0.001
R2583 vdda.n102 vdda.n3 0.001
R2584 vdda.n451 vdda.n4 0.001
C0 vinp vinn 6.92099f
C1 vinp vout 0.91461f
C2 vinp vdda 0.13084f
C3 vout vinn 2.65413f
C4 vdda vinn 0.43281f
C5 vdda vout 1.75926f
C6 w_609_1847# vdda 0.26354f
C7 ibias vssa 20.1072f
C8 vinp vssa 5.42415f
C9 vinn vssa 5.82446f
C10 vout vssa 2.67846f
C11 vdda vssa 5.7514f
C12 w_609_1847# vssa 0.11231f $ **FLOATING
C13 vdda.t23 vssa 0.1072f
C14 vdda.t18 vssa 0.1072f
C15 vdda.t0 vssa 8.26957f
C16 vdda.n459 vssa 0.51766f
C17 vdda.n468 vssa 0.86594f
C18 vdda.n469 vssa 2.0155f
C19 vout.t1 vssa 0.19789f
C20 vout.t2 vssa 0.1781f
C21 vout.n0 vssa 0.82078f
C22 vout.t3 vssa 0.19789f
C23 vout.t0 vssa 0.17811f
C24 vout.n1 vssa 0.57261f
C25 vout.n2 vssa 1.72598f
C26 vout.n3 vssa 0.89068f
C27 vout.t9 vssa 0.30436f
C28 vout.t18 vssa 0.32571f
C29 vout.n4 vssa -0.24134f
C30 vout.t8 vssa 0.32571f
C31 vout.n5 vssa 0.27814f
C32 vout.t7 vssa 0.32571f
C33 vout.n6 vssa 0.46652f
C34 vout.t16 vssa 0.33846f
C35 vout.t5 vssa 0.33883f
C36 vout.n7 vssa 0.27948f
C37 vout.t4 vssa 0.33883f
C38 vout.n8 vssa 0.28863f
C39 vout.t10 vssa 0.33883f
C40 vout.n9 vssa 0.86464f
C41 vout.n10 vssa 0.47736f
C42 vout.t13 vssa 0.30438f
C43 vout.t6 vssa 0.32572f
C44 vout.n11 vssa -0.24136f
C45 vout.t17 vssa 0.32572f
C46 vout.n12 vssa 0.27814f
C47 vout.t15 vssa 0.32572f
C48 vout.n13 vssa 0.44606f
C49 vout.n14 vssa 0.21944f
C50 vout.t12 vssa 0.33846f
C51 vout.t11 vssa 0.33883f
C52 vout.n15 vssa 0.27948f
C53 vout.t14 vssa 0.33883f
C54 vout.n16 vssa 0.28863f
C55 vout.t19 vssa 0.33883f
C56 vout.n17 vssa 0.86464f
C57 vout.n18 vssa 0.29405f
C58 vinn.t9 vssa 0.43961f
C59 vinn.t11 vssa 0.43721f
C60 vinn.n0 vssa 0.15546f
C61 vinn.t2 vssa 0.43721f
C62 vinn.t19 vssa 0.43721f
C63 vinn.t24 vssa 0.43721f
C64 vinn.t16 vssa 0.43721f
C65 vinn.t23 vssa 0.43721f
C66 vinn.t7 vssa 0.43721f
C67 vinn.t15 vssa 0.43767f
C68 vinn.t22 vssa 0.43767f
C69 vinn.t29 vssa 0.43767f
C70 vinn.t8 vssa 0.43767f
C71 vinn.t5 vssa 0.43767f
C72 vinn.t14 vssa 0.43767f
C73 vinn.t12 vssa 0.43767f
C74 vinn.t18 vssa 0.44171f
C75 vinn.n7 vssa 0.24653f
C76 vinn.n8 vssa 0.14488f
C77 vinn.n9 vssa 0.14488f
C78 vinn.n10 vssa 0.14488f
C79 vinn.n11 vssa 0.14488f
C80 vinn.n12 vssa 0.14488f
C81 vinn.n13 vssa 0.48512f
C82 vinn.n14 vssa 0.64269f
C83 vinn.t26 vssa 0.43767f
C84 vinn.t0 vssa 0.43767f
C85 vinn.t4 vssa 0.43767f
C86 vinn.t13 vssa 0.43767f
C87 vinn.t10 vssa 0.43767f
C88 vinn.t27 vssa 0.43767f
C89 vinn.t21 vssa 0.43767f
C90 vinn.t28 vssa 0.44171f
C91 vinn.n15 vssa 0.24653f
C92 vinn.n16 vssa 0.14488f
C93 vinn.n17 vssa 0.14488f
C94 vinn.n18 vssa 0.14488f
C95 vinn.n19 vssa 0.14488f
C96 vinn.n20 vssa 0.14488f
C97 vinn.n21 vssa 0.48512f
C98 vinn.t20 vssa 0.43961f
C99 vinn.t25 vssa 0.43721f
C100 vinn.n22 vssa 0.15546f
C101 vinn.t6 vssa 0.43721f
C102 vinn.t31 vssa 0.43721f
C103 vinn.t3 vssa 0.43721f
C104 vinn.t30 vssa 0.43721f
C105 vinn.t1 vssa 0.43721f
C106 vinn.t17 vssa 0.43721f
C107 vinn.n29 vssa 0.58496f
C108 vinn.n30 vssa 0.42003f
C109 a_610_6649.t0 vssa 0.84459f
C110 a_610_6649.t32 vssa 0.84459f
C111 a_610_6649.t28 vssa 0.88453f
C112 a_610_6649.n0 vssa 0.19391f
C113 a_610_6649.t15 vssa 0.27916f
C114 a_610_6649.t26 vssa 0.2973f
C115 a_610_6649.n3 vssa -0.19426f
C116 a_610_6649.t27 vssa 0.2973f
C117 a_610_6649.n4 vssa 0.25324f
C118 a_610_6649.t20 vssa 0.2973f
C119 a_610_6649.n5 vssa 0.40367f
C120 a_610_6649.t16 vssa 0.28535f
C121 a_610_6649.t17 vssa 0.28603f
C122 a_610_6649.n6 vssa 0.22769f
C123 a_610_6649.t24 vssa 0.28603f
C124 a_610_6649.n7 vssa 0.24425f
C125 a_610_6649.t12 vssa 0.28603f
C126 a_610_6649.n8 vssa 0.75033f
C127 a_610_6649.n9 vssa 0.32936f
C128 a_610_6649.t22 vssa 0.27967f
C129 a_610_6649.t19 vssa 0.29779f
C130 a_610_6649.n10 vssa -0.19337f
C131 a_610_6649.t13 vssa 0.29779f
C132 a_610_6649.n11 vssa 0.25369f
C133 a_610_6649.t14 vssa 0.29779f
C134 a_610_6649.n12 vssa 0.40144f
C135 a_610_6649.n13 vssa 0.19275f
C136 a_610_6649.t23 vssa 0.28535f
C137 a_610_6649.t25 vssa 0.28603f
C138 a_610_6649.n14 vssa 0.22769f
C139 a_610_6649.t18 vssa 0.28603f
C140 a_610_6649.n15 vssa 0.24425f
C141 a_610_6649.t21 vssa 0.28603f
C142 a_610_6649.n16 vssa 0.75033f
C143 a_610_6649.n17 vssa 0.82741f
C144 a_610_6649.n18 vssa 1.16749f
C145 a_610_6649.t5 vssa 0.12354f
C146 a_610_6649.t4 vssa 0.84459f
C147 a_610_6649.t33 vssa 0.84459f
C148 a_610_6649.t29 vssa 0.88453f
C149 a_610_6649.n19 vssa 0.19391f
C150 a_610_6649.t3 vssa 0.12354f
C151 a_610_6649.t9 vssa 0.84459f
C152 a_610_6649.t8 vssa 0.84459f
C153 a_610_6649.t34 vssa 0.88353f
C154 a_610_6649.t30 vssa 0.84459f
C155 a_610_6649.n23 vssa 0.19212f
C156 a_610_6649.t2 vssa 0.84459f
C157 a_610_6649.n27 vssa 0.41061f
C158 a_610_6649.t7 vssa 0.12354f
C159 a_610_6649.t35 vssa 0.88352f
C160 a_610_6649.t31 vssa 0.84459f
C161 a_610_6649.n29 vssa 0.19213f
C162 a_610_6649.t6 vssa 0.84459f
C163 a_610_6649.t11 vssa 0.84459f
C164 a_610_6649.t10 vssa 0.84459f
C165 a_610_6649.n36 vssa 0.44276f
C166 a_610_6649.t1 vssa 0.12354f
C167 vinp.t13 vssa 0.42436f
C168 vinp.t18 vssa 0.42436f
C169 vinp.t24 vssa 0.42436f
C170 vinp.t7 vssa 0.42436f
C171 vinp.t5 vssa 0.42436f
C172 vinp.t14 vssa 0.42436f
C173 vinp.t9 vssa 0.42436f
C174 vinp.t16 vssa 0.42827f
C175 vinp.n0 vssa 0.23903f
C176 vinp.n1 vssa 0.14048f
C177 vinp.n2 vssa 0.14048f
C178 vinp.n3 vssa 0.14048f
C179 vinp.n4 vssa 0.14048f
C180 vinp.n5 vssa 0.14048f
C181 vinp.n6 vssa 0.47036f
C182 vinp.t12 vssa 0.42624f
C183 vinp.t17 vssa 0.4239f
C184 vinp.n7 vssa 0.15074f
C185 vinp.t6 vssa 0.4239f
C186 vinp.t23 vssa 0.4239f
C187 vinp.t30 vssa 0.4239f
C188 vinp.t22 vssa 0.4239f
C189 vinp.t29 vssa 0.4239f
C190 vinp.t11 vssa 0.4239f
C191 vinp.n14 vssa 0.65751f
C192 vinp.t21 vssa 0.42624f
C193 vinp.t28 vssa 0.4239f
C194 vinp.n15 vssa 0.15074f
C195 vinp.t8 vssa 0.4239f
C196 vinp.t1 vssa 0.4239f
C197 vinp.t4 vssa 0.4239f
C198 vinp.t0 vssa 0.4239f
C199 vinp.t3 vssa 0.4239f
C200 vinp.t20 vssa 0.4239f
C201 vinp.t26 vssa 0.42436f
C202 vinp.t31 vssa 0.42436f
C203 vinp.t2 vssa 0.42436f
C204 vinp.t15 vssa 0.42436f
C205 vinp.t10 vssa 0.42436f
C206 vinp.t25 vssa 0.42436f
C207 vinp.t19 vssa 0.42436f
C208 vinp.t27 vssa 0.42827f
C209 vinp.n22 vssa 0.23903f
C210 vinp.n23 vssa 0.14048f
C211 vinp.n24 vssa 0.14048f
C212 vinp.n25 vssa 0.14048f
C213 vinp.n26 vssa 0.14048f
C214 vinp.n27 vssa 0.14048f
C215 vinp.n28 vssa 0.47036f
C216 vinp.n29 vssa 0.71753f
C217 vinp.n30 vssa 0.3488f
C218 w_833_2071.n1 vssa 0.11784f
C219 w_833_2071.t33 vssa 0.38148f
C220 w_833_2071.n5 vssa 0.172f
C221 w_833_2071.n6 vssa 0.24367f
C222 w_833_2071.n8 vssa 0.24367f
C223 w_833_2071.n9 vssa 0.24367f
C224 w_833_2071.n10 vssa 0.11467f
C225 w_833_2071.n14 vssa 0.24367f
C226 w_833_2071.n15 vssa 0.24367f
C227 w_833_2071.n16 vssa 0.24367f
C228 w_833_2071.n18 vssa 0.20067f
C229 w_833_2071.n19 vssa 0.24367f
C230 w_833_2071.n20 vssa 0.24367f
C231 w_833_2071.n21 vssa 0.24367f
C232 w_833_2071.n22 vssa 0.14334f
C233 w_833_2071.n23 vssa 0.24367f
C234 w_833_2071.n25 vssa 0.24367f
C235 w_833_2071.n26 vssa 0.24367f
C236 w_833_2071.n28 vssa 0.215f
C237 w_833_2071.n29 vssa 1.73435f
C238 w_833_2071.n30 vssa 0.24367f
C239 w_833_2071.n31 vssa 0.24367f
C240 w_833_2071.n34 vssa 0.258f
C241 w_833_2071.n35 vssa 0.18634f
C242 w_833_2071.n37 vssa 0.24367f
C243 w_833_2071.n38 vssa 0.24367f
C244 w_833_2071.n41 vssa 0.24367f
C245 w_833_2071.n42 vssa 0.10033f
C246 w_833_2071.n43 vssa 0.24367f
C247 w_833_2071.n44 vssa 0.24367f
C248 w_833_2071.n45 vssa 0.24367f
C249 w_833_2071.n46 vssa 0.15767f
C250 w_833_2071.n47 vssa 0.22934f
C251 w_833_2071.n48 vssa 0.24367f
C252 w_833_2071.n49 vssa 0.24367f
C253 w_833_2071.n50 vssa 0.215f
C254 w_833_2071.n52 vssa 0.24367f
C255 w_833_2071.n53 vssa 0.24367f
C256 w_833_2071.n56 vssa 0.10586f
C257 w_833_2071.n71 vssa 0.38768f
C258 w_833_2071.n88 vssa 0.38768f
C259 w_833_2071.n89 vssa 0.38768f
C260 w_833_2071.n100 vssa 0.19108f
C261 w_833_2071.n131 vssa 0.29762f
C262 w_833_2071.n132 vssa 0.13119f
C263 w_833_2071.n167 vssa 0.29736f
C264 w_833_2071.n168 vssa 0.13119f
C265 w_833_2071.t61 vssa 0.54392f
C266 w_833_2071.n196 vssa 0.38768f
C267 w_833_2071.n258 vssa 0.13574f
C268 w_833_2071.t81 vssa 0.215f
C269 w_833_2071.t18 vssa 0.215f
C270 w_833_2071.n260 vssa 0.20067f
C271 w_833_2071.n261 vssa 0.24367f
C272 w_833_2071.n262 vssa 0.24367f
C273 w_833_2071.n263 vssa 0.24367f
C274 w_833_2071.t27 vssa 0.215f
C275 w_833_2071.n264 vssa 0.129f
C276 w_833_2071.n265 vssa 0.24367f
C277 w_833_2071.n266 vssa 0.24367f
C278 w_833_2071.n267 vssa 0.24367f
C279 w_833_2071.t12 vssa 0.215f
C280 w_833_2071.t0 vssa 0.215f
C281 w_833_2071.n269 vssa 0.215f
C282 w_833_2071.n271 vssa 0.24367f
C283 w_833_2071.n272 vssa 0.24367f
C284 w_833_2071.n273 vssa 0.22934f
C285 w_833_2071.t20 vssa 0.215f
C286 w_833_2071.n274 vssa 0.15767f
C287 w_833_2071.n275 vssa 0.24367f
C288 w_833_2071.n276 vssa 0.24367f
C289 w_833_2071.n277 vssa 0.24367f
C290 w_833_2071.t5 vssa 0.215f
C291 w_833_2071.n278 vssa 0.10033f
C292 w_833_2071.n279 vssa 0.24367f
C293 w_833_2071.n280 vssa 0.24367f
C294 w_833_2071.n281 vssa 0.24367f
C295 w_833_2071.t11 vssa 0.215f
C296 w_833_2071.n282 vssa 0.20067f
C297 w_833_2071.t14 vssa 0.215f
C298 w_833_2071.n284 vssa 0.24367f
C299 w_833_2071.n285 vssa 0.24367f
C300 w_833_2071.n286 vssa 0.24367f
C301 w_833_2071.t2 vssa 0.215f
C302 w_833_2071.n287 vssa 0.11467f
C303 w_833_2071.n288 vssa 0.24367f
C304 w_833_2071.n289 vssa 0.24367f
C305 w_833_2071.n290 vssa 0.24367f
C306 w_833_2071.t23 vssa 0.215f
C307 w_833_2071.n291 vssa 0.172f
C308 w_833_2071.t9 vssa 0.24367f
C309 w_833_2071.n292 vssa 0.24367f
C310 w_833_2071.n293 vssa 0.24367f
C311 w_833_2071.t16 vssa 0.215f
C312 w_833_2071.n294 vssa 0.22934f
C313 w_833_2071.t7 vssa 0.215f
C314 w_833_2071.n296 vssa 0.258f
C315 w_833_2071.n297 vssa 0.24367f
C316 w_833_2071.n298 vssa 0.24367f
C317 w_833_2071.n299 vssa 0.93734f
C318 w_833_2071.t55 vssa 0.54392f
C319 w_833_2071.n321 vssa 0.38768f
C320 w_833_2071.n322 vssa 1.48569f
C321 w_833_2071.n323 vssa 0.38768f
.ends

