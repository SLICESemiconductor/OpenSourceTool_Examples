* Extracted by KLayout with SG13G2 LVS runset on : 31/05/2025 07:06

.SUBCKT inverter vddd vin vssd vout
M$1 vddd vin vout vddd sg13_lv_pmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p
+ PS=1.34u PD=1.34u
M$2 vssd vin vout vssd sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p
+ PS=1.34u PD=1.34u
.ENDS inverter
