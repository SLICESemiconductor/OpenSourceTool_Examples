** sch_path: /home/slice/xschem/tran_noise/tran_noise.sch
**.subckt tran_noise
Vvssa vssa GND 0
Vvdda vdda vssa xvdda ac 1 TRNOISE (0m 0.05u 1.5 0m)
R1 vout vssa {xRes} noisy=1 m=1
R2 vdda vout {xRes} noisy=1 m=1
M2 vload vgate vdda vdda pmosx w=2u l=1u m=2
M4 vdda vgate vgate vdda pmosx w=2u l=1u m=2
I1 vgate vssa 1u
R3 vload vssa {xRes} noisy=1 m=1
Vvdda2 vout_noisy vout 0 ac 1 TRNOISE (1m 0.05u 1.5 1m)
**** begin user architecture code

* default BSIM models
.model nmosx nmos level=54 version=4.8.2
.model pmosx pmos level=54 version=4.8.2

* parameter definition
.param xvdda = 1
.param xRes = 1k

.control

destroy all
save all

* 1. Transient Analysis:
let xtsim = 5u;

   tran 1n $&xtsim
   remzerovec
   write tran_noise_tran1.raw

* 2. Noise Analysis:


let xfmax = 100G;

* Perform noise analysis on resistor divider
noise v(vout) Vvdda dec 10 1 $&xfmax 1

* Perform noise analysis on current mirror into resistor load
*noise v(vload) Vvdda dec 10 1 $&xfmax 1

* plot total integrted noise up to xfmax
print v(onoise_total)

* save integrated noise data
remzerovec
write tran_noise_integrated.raw

* save noise density data
setplot noise1
remzerovec
write tran_noise_density.raw

* ngspice plots (optional)
* plot noise density
* plot onoise_spectrum

* calculate total integrated noise to see if it matches v(onoise_total)
* this is only plotted in ngspice as shown on line 55
let vnoise_op_int = sqrt(integ(onoise_spectrum*onoise_spectrum))
*echo $&vnoise_op_int

* ngspice plots (optional)
* plot integrated noise
* plot vnoise_op_int xlog

* save integrated noise data in ascii format for awk script post-processing
* !Important: Set back to integrated noise data contained in noise2!
setplot noise2
set filetype=ascii
remzerovec
write tran_noise_integrated_ascii.raw

setplot
.endc



**** end user architecture code
**.ends
.GLOBAL GND
.end
